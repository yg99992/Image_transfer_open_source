

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
HJRMA5vkytFTqxtNbuCH60mbf7Is87wQ7cL9WhUaC3K3u6xqGhigYde4mMNOGAAAUsV97XG4mvcT
I7Si6rgTzw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ghD7UoFLMY+hdmZ7V3xXrk9eEbTJD4R4agUb7RaokxaPqc1qoidZ459gXWVCMMkmsI3OlXVolwlc
r1nnwUBrtI7tP+80KOeq2f6nY9N2zDVQaED2WLx9u2i38AX8Yzy/CxUn6BBP0CyxHEePAbq1PqRK
kH88Uat15zu0p+DjWOo=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QFGKtwnLlA8xRIuchvwgSJBkfm7F/OK6NScYKMloBCAApbudhm9TRGDn2FJMU+UbXPCnDGPBd/ll
jex8Ycn9IvFFD4BxNsRiH5fa6kHor6KGTbCnxsPYvEvyA/fvivrd4STpB/WhWyFwfcGPVY8w2++/
keegYcGXcG8Ipxg2EgkzGcIqnpjq60kZX8xBl3jyXLpR4wg7eQVyXgf6qyI9Blpv1ybejt4C3X9f
mWzrJ9+nDQsX7EFJqeZ2ZptWmU/698RqTumsYHWRPx6EjNZdVrCnCwMoUzFLijS/+fY3MI7QQldD
8CLgNYKsSldXjIoGCcoDZ5ZhdAFrZIg3fHF7FA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Sw4139NHt32V3T0vtUGnYNuMPbSXOyHJmtQNlx4+TbSwM4WQ220IFQ6zYuQTg/+mUIv0CuffRVfA
Sx/iTAjq+sdoMdI/BRvTZL092JjbxIuGJwuL7puINMo7a8MWB1T5BHg+RrLTOLXAAEGGA0RxQHyl
Ru1cajP/lO6fEaGmh6Y=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kaZ24FbSwazBQqMgHETs7iZ0cnKJz29HQbRqpChkGN1BtpOIrwMAs2qDjx0zvG6MC4/lFy9dloRk
vOE8g2zisZm3EjiPjTyBee1v2mhFyAWl4xWzHhcomd8rLQImc8G10+eTqluko2+R51AX+3P1Lh7u
+WQx8QhWPTe6s4xo3fBJMPvsdF1lEplAdVrV8kieI7nhdaQPTV3n/EL5d8pRVypk2CgqPyNpVj0k
xQMG/rz6y6kfGp2+dHT/VkNEMGgF4KN3J3+GuV9IU2nE3Um2w26IC+b4Fob+RCqI6eoeI4EMsYhV
reb2rYrjIpGA6Hjq+l6QYY+gyZtzaI8I6Q5qCQ==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
N5SveS0Heso/Xx/bNxrDqH12P3A3WNIUDpgHbX+rOMUkUSCAv9sqJwOg30WPt/hegptCIDnXRcFH
MaEctPQj6XRwtSFggpoLq01kfTHUZBjjCnvb2YH2F7ZPPE6bCtrMRrmPZrH/SzOK/Egy5ek5sBPD
VpDwYTERKHUNurmhpMzPQTD7vPwp0YinzDxvP50XDs4J3PPcWWMc/vpKLwmzboC18Arh2FnVMc34
Qg2A13VktTyRX325eKoZ+dPRdn1q8ZFzMrZSeS2MVT4B0xmVyIs/R3ae0EBo8yfvMZo2mNpDTEax
lhR4gWGlxVcYEMy5jf75Iakyl+WczNfMwrKHXA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 867040)
`protect data_block
gFq+Mj9c0Er+yPbJv67ZYsEDogQR4Goq4YY1rXXvuJ1n4kC0FRsaxdwVXCcjfcGBCxx709tjrTS8
eFmc+GU+VMEcLSTU1gED5ziOgX9JJyXLwMUBs7DzfZK9YGumef9iuLN7NNzCjoHPdNBUtCxYyv3h
ooJRhoWE3JRQs44SY+iEblEU2piFgCaTZDHZSkZ7/fYG7bYJAU0+HAjg1UKKQ0i7yR7La3sEc4eE
jvh7kRHPsk+WiEoIdEE4YgXuD+K/R1fGLJNcY+KG0B8QMCHMYoA3/LHSqLuyRvjdPTGvfaJkJOv+
jH1Hwdzi6u2WZ8fadYf3NY6ZKvmLh55t1LEUhIh8jfKrOsSYkPd9a+cEePmB94HQ2PG2L2d3/H/Y
+/SEtVxvCuDt5/hrG+wNx0cG4/UOGQDJBLGkiGXKld7pjhhA+kXnEMxfuXN6BTERubnc0TBoxxJ4
Tkmp/wOgNFbvP3De+wTYOssgH0YqAo031DupwzE0ncmzvyRlOI60/zNUOYTs4b161A9vTNcA+/O2
FcV84NLpLpiB6Eyj4M8Oeqn2GUJx6+Q0NqFpdGk9Gr8L0CKDSCDcb0yARQISIdQjHNE9v9Ku5MVB
20gScxYjpvW0umNfWGjrnWWGVaNZ3S0zl6Rxy87Ej18SBb1DAsgxOFgJF7gIDZaSnQxRWxXEGX/m
LyZIHTm4MJc2WcwJrS8HeO8mKfBRxtv+dCWwq2xcBgXYe6Q67cJIIXZiJDxSqdNgyhzJIJbxOjK9
XqfmA6aqlVbAnfP8pxLV/pOPEPaY6XgpXiVqygmzBLh3g2chjpJoiekFG9hIyo3W3lyEcz660LuQ
KHFOb98/YhSBLqMs2OCxphbZ2Kvk4tpNHpTSJ0PYfmC/Ruibmqoojbyag5olfW753XkiII9MWlPD
HSpBr51p1nP3tLqdfZoYy17Clg/noIokyaCaiAdU8OwPTyN8plgt8vBINU9cw7EZtAjs5eQP5134
cBjfTTxtsLJ382p+sdDL2XkC1+If07+3DOn1ZnM/dGfZgtTGp+UlJJP+ONiG0wgy55hcA8m8K86X
NFHn1tt8QDabb5o63VobDUFDM30gRf9/1H+f0Ue5I98vIjXP4qM16U9B/ha77FGxHqxwkdZtlGpY
M6zDFSRQEGWfllFhtt2DlrNdRbF9RsAkWW8sR5kP3pkicf176M+J4T8irU/FY5ROz2oXSLDE5HrR
vpLcRBoG9VMIXEbn/EHezhrTHEBxDIa++cMOJF8FjdH83p+7ZNJueyQ4si6NDldNBIh2z5fcerfy
7dq4uQoCSwHs29vGefigZXrylFx1dMWObd64qaL/ZV8zzVU7zg0rkUwlo2ycleuA0Fs0nkRLYuHy
D8qT+/5Gfmww8PjtNYwhvOg+DkUV4HoiD7PiB+W83v4B2QpzqgVjExMv1m2qk4el0N1mMqYtpp+v
196c3n+OAevxd/XpVpXcJ+r63afi3PnztAcDixKKv1OfbKVFC9ZYMDZR4H2aeip1tKOUmLH/+Kdu
H+LxR8T6NMeabmxyT+dDqegCudLZHiR88SMDKPqVcmT6G7OdpkxONDk6TJt1uvutT8KyyYVAhPPS
bMcW/toq8bErKXlykeyDODXEJaAeAsSrmoawURUDjlycwtSzBbkPnoECUFh9Qmah8BKGQn4LKNfo
tZbn/4RyK5GIlyRngvqhFEO7mAQ302Q+1HBfzaHoe/2nogbLsX9xwj/skqMP+etiw7OKKvK2tJB1
YmcsL51PcBVZHL0zWy2jK4tZeKXROykllCLFkSe3uTj5EyY0HdOiGfEkx2c3WVgvowSUZlAGcqIs
XjPcX1+xt/MDgfEL/NLXW/ZgJg9X41twuaR20WKD1PzWGWZ+JEfnEoBE7+Q33QN4ufMc2NRZkWe2
GvTRq7ydjgghVM5qDe/IYWoTawJn7a7BOjfXg3Cd45I5TI3klS/U5trNIrRYz9Zs4zrtnJBxcssD
8u66l3WX8lb9UJOAvg1Z2IJriytkS++qwH8bBObFFMNUr8Hka0QKAYWSF4cM2bOLp8OrM3VXVt8T
HjZ4JdejNdjc0u18XKDVpsPiJC5tSvwiLDZ5Eia0fjuGHDWc2eTV5PX5E/evtjGcG3sdNy+fhQ3e
7FGbNWS88x9jw/ao4OUyciXx6I6EtVelw/7UBn80BmY2S/HKnx4zJvpY0cafXWWEzMivaPuU+CZ2
T3k2LTaW5qBoU829DA/Z3h1jGjEuTX6agVOEO/291ryxRgEGoVna8Nm2nyDtsjIP9PReC7x8CJ/P
L3MxB/eot2sQPED9g+/c42Oaem1/rPGZBrGZNoFH8Pw2cyn+kf+ofIdTux3lmMyz1veBuY9WlQot
ka6RYYC+TgWF2SrTCBlz9Q/59uvomjnTBdE52IU0OUmkcTrrLbqn6l5tUf5fAMU3OmpteJ4KUQgq
QGmmlltH0zxYgkOKVWczfg9v7488icaiIvTVZFAOGCkQwLFjjQ487Fgut//XOgd7QaRns/zVPGz2
NxTGx/aLKBLENqDfEaS3YDHrGR4evi7t//j/hUqZcKLo3Hq4ial6v8J/KVbFN2YNNviEZnA5To1o
OLV1SSmkth/5wRkoLk6hgdlSp8UtpoRfk90OBMjeV/MCr1qcnaYijBvWDAzs9POJ/fm+iYyNv9ci
MluQOPLKJheP2gDNGIYnFNP83fBhsRy0nSQU+/KIT0wMExLzVv5ISUVdcgzoKoabL0NGMi4xGFgV
+WtwtIPi0UL+MVi0g1ZimVdnZ9+C1feGodvihXvNq7K67w9FTpLri8rwrCPix+NcQyQgYfFLAcIU
b7f7765Se5tVM+9Ovrlbs+bV7ffd/nCII3I3iOCxdoxX7GrNyUJQWKtlmphyHLP1pgNDBVKAgL5r
wOwSlcOYNZN8SkjLUSre11fl7MckQE88bpRD+cdJcR1jutZHbI+rVZyMFc7xiQnFvYSsHpJVDOrf
02ebkUsmOrrsg5pTH1zvFBKq5FHKxmB2EK67EdC0ur6CoueXwwUBX1H3TGGCXQtDUbzij4ER0ARR
KZ+uW4STfJ/D/rQ33MOvvjhZ6fO3chM92hkOotNpPIFoqPRo+vzu0tZ+F3zvxQUAplHJ9AX6X4gi
Gnx+nGhFsrvLIR+KWbJnzvtLyWOAIOdXJIw8vinYeKn0ztTKnO0dm9Vve0ZT/h5H4LBNZJxt2T3s
LmWzVl0PXEIVtXuZAJIK7B6cSYh9ql/rvV0TX6cNg5wpHog3gkKNMMYgFm4+njIppu9JWgOnsId6
oNy6fl4l8qdvtCdwm99PCOHf9NtrkY8e0SLWWeAhBcTDW0LysfS8i44wjGOXS7kJoddMInI4HE8I
qW5OVhbVGQryz+nvJdYMAjcPYbdljDZqXTy3d94xCGYHwvVzg5YgwaLXNJAHcv3dRff4Qf/j17XH
7LBS5vbDhXHuhDF46AyeLQ0/tCuJWSaknMIq4LJ8vi5c+C7FQlfOQvY6s8/P8TG8fdtJkKR22sY2
i5r+vjmFKiu2l0Oc6zLs+hAD5QfnrsMOuz3WZZr4I36qS77YEERBEZ43Gnc2OGmXzuhmJN5uwFKC
sKgahVLmCd53Citrwr+SYgcnBjm201EpcuCGA6ERmTP/KZN/Nq6/HdJ/0rIeF7MY49C12mioZ+ew
0Cxd2vNWsTLS7pBwX96HbtgJOj0IFCWiEk+1g9XujHDsX7YEhdVO1R+MJajF1PTM0xMh56Jid73p
n/224nCwo5NmofysVLOnHc8aHNm/TNBKGYoDG1t6A3BzthF9cmWySVeg5VV9Sqv8jgigradCVjsl
ll7PCkU7ZIvLCuwrCEiLZskb8iZormQDG9njzWhAi32eQ0oy5nL4+TccFGEJgOOgx80hv+UNZdl3
PuXlv5BcYads5HdylAMH3TFTTuqPYw3AKJu1qieOrxEdWmbLrVC0hEQthBkuqZORc38MnmuBDuYG
s4slT1OmV5BWj6XqWORYrqILYhNK7FD/s+KjGYg6CJs7IusTcJHFSo+P/unSbqeTSabl9qEujQcr
DogKKMdaTOjLFdHZC6pIfRCGeimN9ISfvZgC7M1rT/c9cU7TNYRO/2NG3GQDE/mMZm9eE+rI3zQN
gLSp+d8hSGFD9MynDnfiWAx7f5ncjJkh+96PHBzA5OD+SPy/2WXRV4Kc0lo6GlujIJRwMuipV0HA
+1ZRU31rTecW3Oe94YRhwPwQ/1FHTowBfKF916OCGruE6a2r/D9xFjdRO2rrPHQ4ZohxrtEVEuV/
DkcwFGx3agXrBn/xow7+uL7lozX4IgfxmI7ImVjc47XzN9VQhDBCDZ6zt3VnGa7HTpZyjaQ+02Uh
8pnueC21KX+EucxutT9oAsWBZh7ovt9TTG6zaGz31pli4DYjpkdiTsOrvcJYEn7nyJI+fVyjsDfK
ftW6Annsi7pR74m02iwGVJg5s2OJ4u6UjKkIdlcWPAMACTeXPJbciZOFuzD5eBH2Ce06xJNOfVMy
kGf4kAwKFrVkhNYHD1ULfoarAmQdBqRE3hKXNTiGP1xjftOi6GrvJkk6mj98sL2+Fqc2YY6pHez2
hNvsr+z79LjLlTt7i+otwhSn+4NyzjpZ3d3OA6Qy6mBD8ErLDpWZBTWBHMtX7Rl4yim9un5t+9A9
vJWZeizPd4iMZoLeoBkLFh4f8w8VpgMMQItoUlRuF47AhvIpJeWrHKH6C7Qwe9O/n8+jzUSs6J4d
ECYm/vCo2lMkv5HVDdwp1slH7EyeQ8R3ImFnhIWmxE2mAvvxM9bjWH4t2pa3YSCj8SpPT0aHvIYU
UPvhIekEUnzg2JF/T0DCv51W9Cuhnh/y9EySin5lU86IoDHg6XzZagnqJdNdcrQk27uxm8/vowrH
OLtcwt/MXXJszGdjDJqqrAgzRxKJWCt+MOe8pAAkl6tX4oli87O097nebkRpgeAgby9uDCswBgdV
lUGsFFawgdPIlj1r0QL9bfA0mj4gNW4P99CzzLt132xvYxgq1op48yAuHA7v2z2rji0bu8aYbVxg
0Y+a5hffao1Rod+CkfH4GUniaz0CPR4c9PFixFDhjuuBazybIDhcH01j8vc0AJS7LaygVtReLbtf
jWM2BOXYvL0ojAtS5wbtGF59GwPpODT/cfckMjCEFdLAioNNc6+O/ZorDmEwHCpnsc8f6weO+MMP
PRxCJBRDjGMa97aL1Smbk+XVY6oitnRNtOplyRnO2ju4AHT5Y2jMKbMj5ZMlI2qv6GrsobEQgQhy
MtQSwbSkDfkxjL2AW3p2DdrZkYkeyYNs8JG57GFbXUE9SjjksF9JmF08FbV/UxylRAHOZmyE0fa7
+vQnjR8EHzSxRA560X3n3JFDVLszGDqQMcQ4xEWRORbfc0rQCLLeWPzER6J84EsYZ0OvNz1gpa6F
wDSuodACganC27EkQe7+BFP6YA43T8H0h/aA3FgJPoXqtQJj+/doRSguxYfMIDPK9VyDsr8xja3b
sRKAsUiAu5QWgVhvjn9P6/6kxqAGwdl6MDDgurjRs68EzSZS4X+6a1D9MOE3LhkOOLLvv/xdemEc
iOVPMDWjyYQuI0yssyFJBlS5860UPws9az4X61jQ8kkp9dqIIIxkyyljculc0lLO1ItFV6/Kmni7
h9wMSP62nABMnYgifLxDpLyL8nIH57mVbRjsmBnMRbZEqjtiyndgzCHtDZlyRUOmsbwWMosqqrMG
inVqTr1frkSeTEkGYmDBwarRt5VawuLgfOlpzi3SxRa6qeWGcAL0eFmj3+Txltua2cAU2HEmOuRG
m4Wp8PwEX9QP24mbE9e64CPT9u99saDvoicEWhU/09GHgMLmAhdIJhvRozMFmRsbRcd41btbDImP
PflsOfQwGCSV/3BGOwzyCC+wpqRAdiobZy0T3DzdJR3TrUwRjzu1be9aAmWC6ekDeXJ2fQVCP0v1
SO80Va9ZjXxndWmRfNcI5YRJJfmnCpPaf1DYBR52/mL2/HTW6epbDZ5/jsA5Q/k/XxZNub2BC60B
v7GOsSUC5KZBkNnaI07WqI9LKDqNFD5ymjnzqDYia4sMNq+kq0lWfBY3mQGcVjShhL5ik7Q1WQEe
PYLTIqBupO4bK7Fxs7HDbmKiom4U1hl7dNDprMHvTuVZaVFmJ/1pyfU6EoanBCZ3erZGzada2s3x
jNEclWQo13nKfUrWc2NjES/IMCtK1gkdhnitmuERZn77nw69Px7y5toYAGUgd9yo7eSacjQz9oSi
f1oNOUy7Yb0plFWThqbsG5L2x8Slx5ySydsPoqrweixmpVfqeJyB0BqJu9errcMyGa5uza1np6Lz
xwTpY4G0fiqTPYi6ZNY9Jo/qXC6UVuTJBElqUuy80mMuMdoxymw5RMLW/cckGd68bLVAuulikY4E
zldZME30BVprm8BwPoct0zrlgo5WmAFZ9gXqgArMrf8TZ5w5jq2D+x2zKiLbURx0HZr3+98npkJ3
r7nlsiCQaEGaOfrTHErtZAFBTn7BNgwTLlCLzBnuAPW2C+Xl4TSVzRf/vg6CF3nOraP32xQ+KbFP
2G/ew9XAjWCdFEqLskOddw/Fauow5Mvt3/ZsVh+cKKXoUbjydT8+Hq7bL8yfqDL3aksXHDsiYn6M
rAqkijN6RtzfeJYbiQ43NIGFGFc/r9HfjBblZRwfStuaHZsX49o4yr8sg4xJu4W3kIkSp1sWDXcR
9uD3WISI18TSO3wPIgU4OL2hOGQB6e+s6dHT/QODeufMj97+7vfsBhk8bEmUHuPisAHHHk7r1W7c
K3yp5Vu0y+YpKGvb9l/7LlmBHpidm/iPX3LAuyvBMPRcNp/PYF8yFA+ePphZW6FJWcPQQf6fMwiA
HIISlWwrxWi+0m+RgKQ8KMq8fanPXcWF1J2xgjS+QohkELmpsOJumqjJOiRdhnEUZrnaYQlLjf7d
yR8o3A3RlAyw4a6NLvLAKCsl361BwbEs92ojN+rJ7BabsYIYiu2Xz1Vo6rvKL7v6BRBO2YrEb9rO
DaRBAhePd9EsoSRRjQmc6XmtjXFjEOS0xzuxV5SPWigOwn7O5wFIS7Qw9Iitg7G3tAjH150/sq4T
Je5STEn+A8I357HvJ50Hp7asCSgw60OHIIVgSXYhN6JxDNRP7naNDBtYeiQ/tChKnuLw2hN38uTL
HKBYqv37Wyf85MTdzaqzExEbNC5Krpjk4L1TCsuc+vxTW4/Czu8OXR9jey627nkRgBystol9oN9G
9pch5knrhOP8uI5OeX28slbpEyNOEt5uSEmmx6OGUiHbo8CaYmdoe0MUM6Qc4GEvJWMqGrMs8XrH
Kyy14mVlJWWiPC8BlVVmIZRT3Lm+KaJVd6lXZTp3sMtVBgZM3DodnvbPhNXd6NUhVntZ6gc2k/UE
dYYA6kjj8hypFCGsGBPpjILUAQB5loO7hOWnGKa1advO9Q0l9SE74LS+Bjis2zU/nFI+OjWAzLkd
BR8/jMLZym3auHDvUHraMV3qQAzKPEq/TTc9tafwi/ghspCuCmss9cIIEL9DF+5lGSN0V2UxUIA6
IQaF3FgGfFpKSla6yN4udYMTXE86FO85qCkLLRLsFem2JkcDXIlbEh5WWw3l/YGLliGV6a1t7rXZ
FCyFgfRlCbZGEhfP1K8SinZ0vtogtK/hffPppI9/PH6iU/wSPWW/5UaNWN1O9oWWLPBV9vhkJYj0
gJUHw0WTUyEbE1jI/ZN9i085blX4JfvrQpapBmBhoyfXuXoU9Zz1evT2uRPwrZ5FcwE59u3seEkF
8cpurVWs81XTCYuRzj6tcmTwMSlb6R/nKjhplhApUPbrHtGglJ7IEdwSM5LKjsOd9r2OyPSZB2vc
434ECWy5HmgAmlPHEli3qtMtO4UtYIPqxkle6XnOpxpzmQ1xuRnEgwAq6gYPFsrO2XG65bNs4a76
uuipCuMxMilzO++RSsrR5xiS+avwVoFt2/Em/EPxngI9z2Ze8BUOlHKvQIXRE0uaBJdpoWkoKlbf
Vqfgp2aC1TZV132CVmixH3qXEOzWd1cbBsGJm2Bvq6iy1Lxn56ydlKknx0PUHlt2bXsoO3u5h1i7
QnTPV6mJjMNxKSDGH8k4LiGiuxzvENgAZhxja2sBWMWPI6idFsEbb0RAXRQXmGInjOFcdStb0X4i
ithmCOzicIprUey9EhCzOQGTCO3veJS7tL/FKqz6sKPVrJys+Y0gZUmAHnM2JXdkoYK48n6migMw
x3uGSrztrArCpSyk+T6VoVB1qYbiiwuIHtTLxT+LihHh0iqmjI2imOpXp+mhSNuMSAhvD8RkEq2s
4yFXAA7H3zZzVPhrGu3eTkITTmPmW4vHVt7UjDgKrfVUpGtWXEqJacbDSE+BMoUeetu0Gw0eis7J
bWZMewd2sDbwUV5+UgGrr8ZlK+TVjrfyKunUnVxBLhprV2iKoJtRgLEWtD4lvT5xB24BpYu7a+42
KY9cRZQOzP9OEyzMIdbk62hwhQE+eu2wPC3u3JZN0wx8UCOdz+F3mFu55pKn30XzKgPTOHX/nJBu
xUFbFAVBCLDoNuqyLiD7J28sn5jlr9EK30z1Qc5Fa67Xeim51GSH3bvOoHNx41CoyPFVk9IxPz5c
pmZLYCx+D58PyTKzA1VSyir6WyXqM2EOlvHPTDvdEa/rCgkcIrOEKOaS+LxxqANWcWJUny0D87iU
3wYEsR1uGKg9dygA4oRh57YWxZFLbCJSrjLbwGK00KnzTusN94Ib6iPDeI7lyArS2gJZ6cRc97tL
GRE77nW4qLYeboEg2Vwhg4vjz7wTL5Nbz6bKm0EI9MWkoiCJe6bLBRrQODur9Ckg66HMAAW+TFJt
/+0W3MxLYD+QhL14z/bj3vBjTjeYe904Qg9cyfF8zJm837kyL62eyuAcLe8YoQcZd9TvMlYpTj2E
iWiFWMnH/lnabcTRKJo3vAEJyMi62oKPZaMc+qx24tiapSWyFIiKFtbnI6kR31rYaWZZJjXeuoLI
3FBOTZqNyiGoM62O0WGHZVTHAsxRC9i8YBEwKX+lbPNTDiKxDyrFS5x/sFEew/NeJCcK+i+t2hdM
h5PzzS/UaDEDp+QjFi8jJvYuayZrH0yJZMYTKRqLT46VrbuZk2bhdBW7lz4Wa5+y1nNHateNNkWV
wrd8JY4SPIQipZximGRU3NQAfwo7vPbjZvcvg4Y13rrpb/Y6/5MmuOvUl1pVHBJkeHvjaNA45myU
A+Ou+tjf+xl2/xWF+7H+A4biEnJNNpnqYg7Bkhu/HS2qL0cMrSB6WetH0Dj/lBPuvF7oQsakhThB
/5ysa3n+aj9YtVBBMXtnd+1j+U/D4fNSvxsU8Ta/legKDTv7lDcYA/vjYFMQrG+MJNe5M0pRMsBE
acVGj/KBHSkDfb3rxPydwjYIoT+pPfZB9NsEhfOddgCpuaraR7r7Y0L72dC/sJ3bBliNvMtOFXPt
kTl0kbuF7e8poFp5w6dI6JeIEGI0FBcCdRag1B2/EblZlCqtgn6K7xFN0ioNr2g2ZqHBPhJ3LSXB
Bx1rU+oHmoXtLrYnlHqwgwTir94/Yx2t1zSWlFHo4OMqKg2NgfkOPt3Bv/GfvreIvYc0CmTNHjnv
g9znUyH8gVcwdx1mzNKpbwg/E7zDFUq/RjZXldAfX63ZQsKRa04pbzAmc3ohNTqQdyAiiTWe6Tbc
ASwEtk5aKK9HUYxQdi6inoVFvAwh1iSD4K46X/TEUmFNympJ/QfcOCcJn0/kdWoXvmEcG4Hvn7oP
SDgKbzooN6fv2mJmSnrMFLqE+QxmllOMJvj3KOjnzsgp2m6MptinTkH6kgcPVNGhx5Tbl3EEzSAh
1smPYT5hj6PHZQPmNO8WMtcq3AB3M3cP7vhsubeUevRyApTt69QHYBbvDhqZNeHToRF0hCBOwWOW
iZszpfSAyurwxkI4MMaD5XEPLq67cGzi7MVXCurGWl/n22UmoznmJYLWYoAjqRIYGZzaNm6zbnCy
MPcgVq4Ks4umy6J1SUvYf1y5WcurKi4ROCNgRAIABaaLxcDwmUq1lcFE3U201VMfXHcF62C/j1UZ
pKzcxJo5q+SyXVjxw9uWXS/nq7LFth/QSJ5Jd6uekZV3prLKka9LAmMXUsMrt9Ba3BJJDV08RynQ
Ys9tMx/lC2ytv7TuUFaZPhitfqrIe/5oV8ml/lOPr43tlY4CDk8GZeWbb6Xt2vH7j9c2J74TzLkj
6+s9rQdCsVEXBwTxsVrvJYtz3MruajFwK/qPPXaQLR6tpQzGEdMi8KaEWIt52js8bCik4fELktT6
fu96rMkKviD9x2WrL1fO1fgb5VGF9V61jXMVyb1SJGcbjuhwOcvrL84s7jJ1Xy+hK8I1nGZ0u1GG
nqVYhQPiPohSgQhkTmILSXJWf/Q0KOUdUZTb5NF/sUkf7LJQT4RWjFUxN1ucIMddSsmXiiI4Ov+Y
q09XSxKhv3wid7G9ZYhXgAE+q/pYudnDA2giWp5mMSo5Hh8ncUpPbJqxnuS4N8YPMKKDgUCcTRHv
VGcRQ2KoPAr2r0rMw3ri4ST7t5dycs8S084x8JOqpvl23GuCja5wOua1xkQvL61rK6w3py4Poh6f
3qxgFjowBuCe/Fwk24S9RD8BtGNqlMuhl26y2ZVUz31xq28AKEh/rNY1caksEh2ODIwnAguqqio3
1hbCA9FnxwxR2eQjd+6gLxETUQ4SJN8ChOacrZ1WO84HpFv9GiMXF+qqFJJYu4MIjFTjABOJc5EX
AJ0CqpODodqvRTftBUvTxc5o3aAFRGEvJVa01gLwXM55C1WQJlGtgfn+/UZ39bLnpeXRI0WHfmkE
UnTgRmsq0IVyEmFqWoRnJuCyKHA7bWT7pvE45RK3mWl3W6EWzGOmkutc7J3YyOdYxsGvK55JsvgC
ugVkKXHEc4pUGNaXzV8fU8hO6/FJjSWEn13RTShFCYyVOXn3MjFYfUv6qUVyctLUzO7vvFu8fA0j
DCsJS1kAfYfZWvFvh4LAgMr9tT1+gJQAvkmcl760Fu4OzJ/fiO8evAorJfZQcagxf5vNzEcv6dbF
9vrMpee7l7nJHuEDqXlGbiD2vWsol4JSfhgn82SRNno7BzeYeESvZcnN6wcj5XCduhFiyZteriT9
T+x5CoINnElQ0jXWccRGFoP1Fs9kV87NGhw3WulRCqUvogTJjodm2bgyL1W1KuXmfr0nwgCy8Vvm
qt/ftriiMLk1byA7HRbdeiMPn+fDNfj7F1U4z/3VMBDH09dEBIb1GLR6y/Jc07lmzTq8ShW+5INl
331mOZGUFedBLqUHf1GvntXoR+zlgbp4Cv3TvQ0I2KsN5NtIVFd8F3rxJxMQ1ZnATogX8eWEMV49
jm3kRHuzDhapYiO6hIoMXcOstiYRWi33o6WivcJQNrrX7ueuCpUxvxWcQATUhiiFenB0CNIJdn8W
xojwPKDP6irp0eS6HM6lVxy9RQOuagQTif8SZ0HDCdL9/Vo1+pB6D1X87RfL2v8iDASim1FDKvLC
E3UMBZ8tH6lszoCs9uzBw4LfJ0VUpM/gXJJrxTpfNwwr84kdtSmrgsmRrBNAg8j/K3FhC9ZC7Za5
kN2DC5jQt0U+33CJEBnwzoIvEhTE2cY4AlTBfDNene/nW0UJc1LmTrBkz6AHblb7nsGJC/DtgZ84
Hy08c/3m7RF2Win7RHMobE3ukxentV3Q8DLs9S5dj9dy+PSctRmIja78mt9Zg4Rb6WKgGwG2MsvO
3P3Wh6ZvuShc4tsfjuqVlU9sL3IXAxbJpMYC2VMaAdeLxKe5qTeP48iJJdQAYlzOpJJ2Ed2oQbe1
ZT0aA8VUrk8JY1hzHypJzDSx6g37cQ6TpwwmssviH3EnYev7smCwANNYM/O8nk0KqSVq/YEzl4G5
iT8pNEDDbP7vW8rkbDwkvtE1+T0U6XCsg1qcvNX+ohgjGuS6PJEhdVqWN0TXLU7JZVElbzZnlkRN
phsCAxJLTvb0oWc3m9q0z81RGgz249ZlA9kLWXf0ZPVxR3370R0dnKUKhnhC6W5GqQczjIYtWmKj
Jg/W4L9zyiSsFHsQ+zx1TLcBnfezGir49A5oXK8+R6Waezh51/yKSgk/fNImyIuRqC4dx4IaLg99
Vip2MeQRkcXh1Q+dL9RU4oV7HK9sSJvM8RAnIi7yjOSEJmrmr1jRWOCzoso+BlFFSV6DX4hr+xEO
DZpEXk1vMwCzKWLukGLYsLUfjrP9c5BdIbo3WShn2V6ifYmO7Q7naHl1+3iqVblww8XVqq+WEIsB
QMJ/7eOHTgzIZ0yZySXxi1rL+Bvl5MmD83vscDen3YNQf+UAEmKzt73Vm1gLvwub+2HsukbE/RGT
X3xPHJazsYFtaC3mFFJJ9fznkNjkj0sEB6s7mas/tSxhwfa/3HS/LDnnYUn7H3+pbASWVpplmrWe
OYbWj228QyWIGlMVz+B2u8hMqVK7SdC0yndHdZvbg4dXdf4WazY9BTRvmfzBd00VbnTWpEsmq27Y
Cd72BNDwvMMB1G+zXgEVIHcfDiGB3xVfAabE2l2DJi3y/Id2/UO01YiBdX5e+TDv6xW87OL9Ka/b
S8BOtKkYLA8VznZqpeWv4QjTvGEpVqt2Vglu+O40sWPYV0F4q2l4QtwwFqQUa0aP9R0l11+q/gaE
WOrqK+ZUH+DcTq1b6o1IWveBXcuQZ2bl6ceYz0L4psi1Z4VHnDHv/4kKOGpiJQhcxkYKhfCWXyE9
Fgo8bjPlC+MqByZo/B7djeuD57kQqdiY9jErvkEbJf9R9AyH3cCNh3FJVJCTt0momBDPFoPEynpL
F+IK3Yma69InncAx0u0i+UAJtUTH9FfwwqOxCqRP+MIUBae/WREIL33xQW6q4L5OGFXPsH/xtVVS
sHBWzJp8fK6ARMQ+ZO5ALGW8LZMvRU3KrhsVmZkFIvrAdSjpcMmYfTYeLqEmOA8obZu0/XxY/FpC
J/5FGQ/QmfjUeHYH9//u1VkAfuMSqT+rhFl2yvYVkTk8qxJaN+FxG92n1RGYWDpJMMlzsm8Y/5TD
+XLlXKQwVmcaFb4oUYFKwX1Reta21/84gKRv/1vuyWzxxWK2XTbSFtV9COr57f2P+w8iWWSbFu6B
8l8wD5kzuGHh+/GfiTMqGyGYOy48QZrGkbOwW+04FPdze3diEHjQaRHe1R0QNI8v/eVSSdCcJc/O
IRhBWkovxe5aTjhRP7aCu6oZWskIN+bn4eGzLDMOj1KJW2JWGR+VyYPWh21Y3G6CfKVX1aJuLX/b
R7Ys0QrsxAFVthwKZn0iTzOWi5MgNBlDaRW3v1jvxJiAZOB5zFlHoTy+cTzgnP8YhAxfXSScFtZM
c8ZFlBQBfSKbRZ7bBJGQwj4gQyVm6d3kLuC7QpIzihoe0XkPJmxFjMcG9akt8HixFYaIItMjejOC
dinruHAI67kHCgUUlyj8DMzBU1ORYisuaeGK7Q9nHGpBc/Pk1ySAbgclch87+dWPMHguauJs1olR
0ANneedy6mbWqBd/eGqYjXAU70Nq7XYbvAbLboZ/N0UkYCib69mmkvDE4i5iWiP5qYfV6SsXj7ld
MRg8kFHczUqCSnWQK+EIRVInBdo/84j77iV3JevPynx8dFfwz/9KRb1FpJWSZI1s0O5/uZ7KqEvM
6X9pJ+gt4W4xei7ovMPgTlJwXOdujKlKYyBeFcyU9ItYw2DvvNno0RsrHgGgIrTEJhatag7V19ln
6CiFtvXJrEyd1wo1fIIcv/PwUHGiBWqMixG883cDXUBgN6v/8zb4K4nfwZW/gsi1F3M22HAmKMG+
KHYsh9OfW4edcrVHGnOGHsY3wWfm0qFpZwMv7J7cZPEglpBNAFlVgmwUyByMx1xttDtq13kbhN2v
zaUBVInnNqcoksdsjuRWdxWrPHRBXHYG6RRGwaY2v2yS98UZNNo8lViH0zLZ0uedfnFUirTKx9KF
YrUGB2AdktcOwWeLkgPbdPVlxWuXOM5PpnEhwGWPeJv9/KZlnsm2irzNbURQDDnuTSh7RDAc491R
bjiEQogDgEFE4noC2yA3BYW7vQQoQNtr1I+A9VWUn2U5tmbVQnZm3D3bYt8CmhPUvPojm4pWGFkI
Bz/vcHTusBOjgGlT1U2tirXW6vZS00R3HgeHqgmca3V922vIhRjs42gXEOJv8Z41g6f9RoGoiHWS
RGdRlv3nKIihCr/00EnG4PgsWaUHgs1RO06D4KvXHVHIsJfLGlyfBu4j9LhqHQGQzRhG5UDkAcU4
P6FP+2PWuggCQIAp9b51+f/r7soRNNiy/LBZlo7oHem3HxjIP/K+xq+qxmPDfJgpL59/kwUBjCRD
yPsqhDFt4UfOoM6cR1ttEd9N56uIqPPWetgaXaP6c53V+/O7iF96mc7fM9NeasK1foLSC17W4G57
+v/zFr+v+b9wI67n/SbCbU1wGf/XOwV7uoJt7hnt8upRf9VanFl/2BEti9MfeC8WK9uCNuYvQo7E
RQW3f2q/zlC49EJonXX6A53wnh8K0UrcMaqJpKDWpoZwGvjXJjmTe4e6WBfC1up2kcwv7G681O1F
pQwSvEJIfzGjzdn3LiUijz947MieyVMX51CD0VkVDd7zUKo71C+BuupUIb0YaSCm3fl/U4j8wnFF
YYiJeARq5LALK0xoZX/uYwpLE2YsyMQIVCE+W6d9azqPv4iCO6T1qtnH5NkUM65DQDB4WsF99/K2
ohDNFMXCE+wbTpWM/rTh+IszOpp1wHaXY9ohjBVEnliX3lsOedU8x+cVNqw62b4WE/8CbrhT6p4/
ohU5gNkPkEcuLO2rqESvqFfGu6mmjgsq4sq4RvRzgzuUdZkjd8HRMzlWOK8y1ypYGQ1UnTI9Bm/2
ov+uWGhBPw8weQHfGJOvWPn+BazdkXFvM4bAnrL72m5yoh9zWVKORa9QP11189L6+u49wp+yelsm
U1vM5ZVXbzzV+WSc5au8O4rnPTC7TdgUui3W9YYe4Vw9Zvqc34Ge4Rrp5Tj/4Ihhp1CBHNQKjRu7
JwDfesnN3r4B9GOWL47UimDnqUJndudLlrjrw9/CB2i3afgxCEvuO0gTlFHJKAIxFM8jFsxey8e6
XzVpuhjIXvT9MBygwdyNTRyjAG5KfV5oa6d7wMBnkbjN1q5Qbc1mJwVzSWeJWqzFNLmrpBJM29/A
8nufBUBTo0DS7ZvyZVIi7TeJOzCutLV2qra4OefL+iRCUwEwT755tAacmQMo3b0Lo4Us5HkE8cTz
g83U36tQKkQEx+lrMDH36FauvHG+/hQag3dJGyz1kn9bHhSbJU7zTyP9Gb2Kq2cidOS9nSDYQ1Wr
lhlJOiCGpbQgm1DsFkYP+0POtlSS9wOUkSPx8B7F3spHsS9oxb2jCgmMjTPhRkNG4LKV/JXnPh8k
c5ytuhiiPFqmdQh7DcPaC4kRUMY+evSijy7Ky+UyqJ8uSs5uSP5+Hnl+t4ZqCuQbr7Pfp/642mxe
U1rVeRTmxM4rptBNTpOpyL+wcOImFP6pRPpgdFHjpeTdsf2vP3TFJCjzTQLY0F+LoCGBfqIz3MiO
DIW7tL1xa/X5dP0b6LPqfp3eGMNPLU8uxqokfDLNMWo0PH1VxP68kV+7axmx/x2AdNUGBXmP4Ke2
ERytc1k0HOnTDWRzbCt2czzYgxljMiEC4WrqE2AhAFWUuGTzFgLtzRWT0LMkwm5fB4StC4S+o2oF
GiusnQFlTyFZe1uSzArxfIbMDeRyczFb2/foK2KFt1TnyralijTsH7dilWqDRLVecSaK3rCjlt8T
OjNxXjFmynRFw0vNcnf/vLna1/NgOraaviI8MrFwbfMucakRt+fbYzJ9vjhXZX+uGrQo01jp1mR3
RPBNYOWFiCPCUg68qkwCqLx0Nta98qqwzBobh0JH2LxJMPxNik6XTFpo3T9QbTd5Av5MlSbZa7M/
wjX/OkcdDVG2vMjzTd6MOMPoZjk87pilDAceVzEdJRkSSTG71x9D0YMHxwYlZaxZtCYix27fvqRS
P0ZIu6LNwgwlZbcoDgMdGWJLOngsux4Sm6xpqOuNmkuII/Js9CBuVe1xzYj5yA2mWXWAPm7eDnNH
pahxzkwwiEr0KjHlVCzwL+vb0ykH1sWwTY4cTxezOluGh63WQ6oJqriGwD7pcIafL9znZI3aWEjU
+Gf6nzZV6E7+r4iE+MYERY+pKoDZ3tYJ3pCWblAaZFoi819Nzxv1lpdHNlktWwvPbIjxmvSoitJi
LPJM1MGqMMmkUXahAHmyFWCcyPcDYWWBKpk/6HBmGw8rcqccaHeFPKKf3e2pKgIxO+pk7ovSMdf5
3GEbMqHbAJdLeHWAaU4Myo6ao0LB4auhBr8EhI48BbL5m6/EX3VV4PCUXQGChIPX4i+YRqZVJNK1
Wu/2UHgyfQB0pBvrhBsPsmv7tYIXo1WyUrcUy3/OT9/zBAQOq7rWlNwJMxaFu5Nace4HSOFM37G2
QqMiHIu/aj24EkmM8yvltjDn4iq7sAyE8Pz0kRezT3IO4gRiSZ71rc7hPep67P0FqpOBslsCSwda
ZU0uJoI7i7mB7V0UibNW2Wy8ybxHVzxvbgZkD/gZwgDqw+dty3uaDGdWCDezNxxwYOYjOgsgsQ7r
SXGPS+gEslx2eB9+A/7Bk+Uo/acal6NSXy/X32rQjK7hOX78mfBRCes8ryCHwg3d4HrK6XMtyHnF
qq9l4QaaT5mwXiLgdoFjrAnttoy2xpYYR2Z42m+lUvvWMqv9RcFkG6N0U42W75RhaQ1hw06g0TFY
kscZBaUGz6inhLegYUbxUhtyqL9swB7IIHEIgrv0FSTQzSLSKEydB92KIWv3/wxKOza579qEUhKY
ZpnrhWJTB5grnB7FAi+876jYpvLhV2OS6FcXbaP5lHPvpAtvIYHYCnyXhj9uGeTQsHyqddyZbXsM
Tthgi33NqsXnDr5YH01Dv8mz96rrNrrHTxTO9EnW/ndsxpap0gUZnsFisK0EJzQDDVv3fCMBgQ4f
mYQSru9CEtYzTw7RUigeRo/WS/1MM8sJber9Vd9gPwntykOtlDiJ0p1/M5VxYkZT7t4ewCd1JeLI
e6QMGIgB8JOsLpmOnHFjodiaczclpPzGXNkCtJFmF52orVKF7tEONvnvHs2UtfHBiKXRkIbCUXL8
EBc6I62PSy+MM7NuZ2KqE+AI9Qp6yYubtgNE4w2MwQJjFhgiLO+OlkBPdwgQvik33X5iqNzdc/UH
TFG5jIm83GZf8NUBtuPdR5vGacZlEF6CIjfZVntphBukSPXuDqNLDwfGxMjvyXvKCD7fvp64vKhw
vsmcEQXpZrvdRVZ3xK7n0zx70ORAIW1GCS2JMEA5PApY5z43ou35X1m6OJ9De0cnMOER2vJk+bEJ
sDn/WL5tn+1kfyhtWHy20hRIXxiKg/JKZ2zLohdgPwGL0EVlpHMOKO5nwUlPfOF9Oqwy9XD7qMXD
tlmntiHhgrDsrTnhEQm1mSiII3DfD76L+UWRbEVQIjRnpXVmkxAEZ1HT/lQc2s0ArwdyAzCUgIRA
x8rRuiUNYUIjTwQAWdexK2yImVocVoUFZfqu1f31AmFaJaYv8DtJPwyhHTNlEpEdxgSSJEIrP7NB
u/pEfgZBr9w2cyPjWjeUTHL7DxLYEby6v8a0oSg0i5c2JTmu/zfICaXTbIB84UyhMR8Wrq5TEjt/
T2DHlJb8ZR2CtnxThcbS/vbziHqhc/wjAEv9sy9x4YAQwsuhiLD/YA9CJSw/jSFV/m3bIhH9H4nX
Dta50v7pLtYy4TxvOSrQmbE4z2SvOFiYZMtQP7qSXTBHs3k2SGzPlF7Pxp/ToNDB7gmN2Kxw7Qme
4RPFC9dgadYvaM3LKpXS3shUPfT1tWR46JF/DEQiRUoQplxmv/2lI3MqUzuKtEXOmyMTOipHMwSW
5BQ03fUvEMsOq42rRvnGA5tBgp9ZTvmJSVoTo5t6p/xcEsjpOT3LHEacUv1Ibkmg+DWxhEssaBwd
K5e4HcgGOE89IuxzfCq3CLiS517Cp7df11XlUkTH/3622xIEOl6OjjbSPdFeD+DMmGLH77T3FmFf
lC5syvx12wXyo6B3Qxa1lIbp5PjkQMh5i3aeQOzoQUGAv65hIx+9nQbCFvFeIArNZ+SG1jt1oUW9
htIk1GQEa61YXg91mc4ZBOzn2H4GYywsAXvSqDUSfo7PJjlibn9sQs0KWgAvah1lk3+hPxeV0MFV
O0+6Pqpdn2Xq1kJra30LTmMNEvfsigplxlUYC4ozv+wF/pCCT2y8eq8oyHJdTsJtXg7NDAv+akT4
CmUuKEFk9r2acXlt1tsBk86xNX2/wWEBtk0Jo/yoho9aRNFHe/UDTrN0UfJJPiaHMDlMDKDdbDCT
RcHoaaJHO94x+rU2f5eqwwBpWD8qwkPLs9srOBqoGxM+3tShQp5h2/6qOA3s9lUVdwT3YnY9+WzF
Jup54BBO/EZ2f8SRv1nJZEhXrActuxfSsjvRBNRD6bR+vYvCwKVnjflkER76Qq6LnFyd3GwXKlsd
ReFZaPvqjpWUch5qMRKpRbw06EUvajNo7fJxIocXX+R7ZsmoqOEwEm+hSmgBL2ubApaYNJH+IUcs
dBwiwLnMWj5IBL16inoV/BwZBtEo1xhLvm/wrErIjE9OzO1ccDkC69uaCHVY3aOda39UxpcouLPm
9whTWVLfFYZ8tiu+ryGIVz9RhRb5xKFZio17/Mi+YTpfskhTb0KiUttCMdPLfRprTePONjQzOX7A
l6XMLfxJ0hIj7GnL7B67jKv4yt2wnVQ8GfboKi41Seksj0fL3XPPdbhYvRyi0cpMqClPwnFtydU9
SFdllZTG1AqLN2ItnAtsHjg9lpsgR1FIWAOGACjeKa/gmk/Yv/IYFRyz/lY9rZS1JYuhR3SiR0lZ
GHVpt951nbl+FKs8pi5CvAdWy7pVRVE/gICiNjy1hiFlMev/CSpqDp1eLVtXxDBEJf4DbHQupUHJ
m/jFVuIeEs/2JAKwcV5wjkEsjtcD8XjKhbtvL19pkc8zoC+nL5Y+Fxo2iWrZXqSlACXpO0EsBI3S
0kNDwfyU5L8Kj0FdoR/2+RaUymwHnqYfin4QCqJqF6GwiKf5byHPicGZV76Olpdqnb7vwF182FPX
s8f3xvECI2XzURBBJYHlwh+JuiUEDVdo/G9opKQglEyN9omDBhYTrGpQz8FHZU29Yn/bgO6WGJzS
iWlsuCr2FsabYsBd9hVtE6I+L1g5tKqH99EwFvatQR3TrC2z7Mt1fePkRpMqoqkLmDyb6zyZ6OnJ
faAc5EMmF6XZCQIcreZa2jC/sV1K+w5ww9AxcBkdapTI9CNQs8qlak7IYkOWkQyiZfsNOFWHRpSk
0kCowDPoLwgxbf9DqLTUy+SX7vaap0XNgDeBVI5pgsnvItvL/1k5zdMlcJ+VqPNE6kFRASVWzSXb
hxvTpz6hZ8DRlioZDjwHZEy8UZXkV4JGvCWNIcphySALI8MKI6l9LV+gc3fmN7xgOcujmVFXL1m8
/iMRGJPLoQRpu2cE11t6nZgCRzu03i0aVvfStmddgxI4iGWxP0Qbpc5tK6Mvcd6E6FO7HSRFCQvR
fA/Mqhewv54RXm6FmI0pTkv+nGbjYFlhXTtyCgxrg4fOFsK7hNWRxdkAfePDepLdnNxwo8Sw7i9R
9YjVJBatZgNuGEVBHCkBcSA/QlTUVTOy9m9qkG8iQ3CbkwIobaZ/mp3yxKhi7NZU4+3XgGm8NDtZ
ZVQSxMqJrgWFR/RigzrpQG3mT3LjPODTYU2z89ccbU4R03JWSrX0+f49w2V0pDCZIx/i1nIdKGYP
iR3uz8zO7UjwfGXVjP8oSrtBJoxq6vmM9QjgRXWcaxj2HfHOj/K2T863Q6jyuJyeoPUVt1rc3K7F
ISBoaYz7ycZpVC0KmU+PebPXY7xgukHHVSlH7mRMm1w6nXk2+lVHoxCj4NpSKRXjtE0sDC4XEGf0
614K9D/RnA26pJ1j62+iukfQ9pMt21mPa2bAEVVFk5/CiohW8jb0jQYrGboFc76QVQ8jLNpbkNU7
0TL26/IUrjFo8wviOv62KIaFcCZm+QcEzc/la6xL5682Vte7H4JcOVwAR9IASOxDFZ3XKY+TVELP
vdhfvISSJrW3h09Xs/KFrtvn4lyD5s/0XmRRfv0RriR7FYr3qPMerUGgO8gYiLOSvvY4uCskl0xr
xPYQI/SwAYt1P4tDPZ/mJR99Te1uDRMT/vYhHFHCjnCW1g9q/+6YE5PniDBAwvS+aHimdfiBsJx1
B+FJDg6n6yMdLVATEyYZoCB1qz8Rf13l8spaGzvAxysceJrQjvYGsQg54rLqBuMk7QHfHZVCp8Zy
enT7+p29NiyXjaid7wn45LQG3je3M4HXYP2ylOA3zBVpb8qUUfjccZUheWhsviSbEfXAJ5tsFjKJ
I+c5FPT9fi0JEp4W4LGfGRYPHlNTpBTe+YMlaTAX+0Zm2+4IaOx8CJky49ccIoGytQ1zCtFtBfYI
Rtn7Qm5PDEzXqypduaF2BBaaJEQYvnDjPyycELcPZf1EvYAPEWAufB+wok5+/D2EhjowV+KdA4Cw
lStOB/ef8tfzthouZuiGfZiKjyO0pknZVFc84J+AWlupqR5XyQ9LcpfuR3DyuxpXGr3Zo1HlPuvW
7+exNx4zloQ3JRVBBFb6sBJC2ka49g/OIvDJ5Fz+qwFj2xyHvHv6wCJx/JuhMrC+3aCXcovgQcY9
P5d1gds+w76raNvWgyueyfu6uvCpOjkKLaLW+UC3iW26gK+aPvNLHZFDKn03hlTttydiAcyXL5Yq
kt7ccH+VphoTnY4YgOOSETXoMb9Qg9PTa7dlmCBLQEXog6ohnWh/BWhM04nu03tbp9pQygFdHh5+
CLizL2+sG81kyian1oyurCEgbdogsPh8UChj8o9RIzBqvBjo8w4JcmVshMvupHxt3NbrAPw6j2HZ
OB4YYn4zdgjTo9pQFzKVyuHbxBbBhmnXOc3pGxIsjMcAkfYlGokMPOuiVVSjyLLYWsZb0Qmm5MOU
Tkdau7jZRLh7Q7+Lyc7unlnn2gGuT8DQYq9jY+HR4JAZ0B+hivc8sUiTznOIL88AuupLvayggJnn
/Z/ULF39BOJyE54Q1Bu1CXPNnPbOVZAMirfpwQ9veCJT4s44FUZrFet8CRtXQP7FIREgFHdS4HB1
u8mLRo69kXXSTXwUFW1ZNvzj86YvqtDPysEKE4U6jk8QME/wrCCQA6v0dsgCrcmuqdQoSAve3g4u
D43DFfybW4Wy0Mza0hG2aQNSnb5Vbin28K+ez9KNKO1SOc3ZJ+z0p2ZuXV09zCbvcvuBYxSihPMR
UBAS/ZFawLEVClpRfqYf/RoPdm0W59GaaZSXzy+AeZubx21Ozaq0fjsKg9wRAABnTPtzedDaGo42
wqTxlYswQwtaThcVABhiLh1cOJ5v6UcwcwHTCbXNWNcWuErOKJ+Prt2OYx12XhIFL+8XTmNU/pwz
j07oVfRiUANrtNg6s5M6V+HhvzHlIYPsOTlUEIpZLIsPoO6vTiONOndKtGct3CQQNY7OPXjzdPBy
Mk5pqdPle/+odBofb3sYV3va1OFW/gB/znoGd24nzBq6CUjI96Kzmtn3es9IbdPEpd25XV7++SWL
3BAEJwU4EiDwfNumY8Q+iboZF/1lgHOKULJRw0qjliUx2kYW9lP/JLVcvZvAusvmHUs8hUopYqdX
YZSia1JLf21CFCGPbgallHVFw8IO0FXswhQpl4gDbJdVUfJ7NwMx8JNogoUo64JY6+v9PC0g7tHI
BfMdosqAhVPUW+sExvB125gvIxEIvICMwhCwXpxC6EC1pq3dbhMahPiyaAS+OfizgrF2OSIyp5UI
Vxauav6Ms3jqQHdfdocUUhtlT7G9WixHv7DLTXl0SWf1uM5EkndNiFtncCsVxuqSSb/vJsuSYJU2
SfilytfdK0olNp2tohHo3JPBYcY07vfBI8gzONAnxs5sdxJpRcClV0le4od5BcuyXNsW6F7Agm8g
qO/oDmqFR1BTTPLBb7wEK1uq/o9lqpEhI1iuyiSz605RtPFBcr0vUOLhYO59mrMIJ8mSe6rINsGi
jkfYFeQiA+enHPyXOcwopAbSg6z81hYZqtnUMaedY+pL2rNvvzPY9eU89G7A5R/Arc5RhWyo9Edl
kyzQlYaAZUpc9D2VdA42b0+I8R2FpE90IFI3mXQJWXzlS1v9141pndYlwBPk5dHNluQMgJAm6bWE
aKwh3RXanbpltQ08ksOA3drJcnA/ix/YycEH2h+/IB30mVw/P55om1IBL2b3nNsjpXEnfUAxS2fs
UpYql2EDooXTVeKm8GXyx9t0GzqGWVc0jzljUfDDafy5EaLn5rt5tna2TIhzCdVzIycoaeqGMziF
DK/RegrWU0bif9boaijtVKpGsLREoGnq4aFhgPspIsm4m6/2XankbAxSqxALAj5T82LKQCn1VLzh
dmIyEeXFohhTXra4CFNfdBlbtvuXBruEL40rDmWCnoFAClLU78TrKEtf3j0STFXnRp//N5kPIrfJ
ll6P7Zgjm+iUa7bsh9pdIPnIhVT0TBal5Wnszh2K1EpxzlcaaubpaqfCnpfEoi12n4mcRvSPYfIW
2x76SjD/eEu3oiQ40JCwUO3NMRr5ZvEsbPPWbdu7Gj6FfTYw+xdX+0zxbkGJIZc372a22pHL0uAM
Svgo5op+Sx5YYL2vEKnPTujXSNR2VcSyAX9GnlOYiwgPnFU9alYzjNyNYE71/APIn3MpTFqiDxyR
Rj4qQWGEs4qJbB+/+Q54bHTykVEOZaWPkBXqqWjlwIWf/9xm0Sq3En9Bxta14Ge+jnYpNSNkkv4X
RGhycIgHK+AQ+wVyakl93ZoYHOaMu3dMT24sNGzg4aO2eAGKjXZWCK9ACEOpuFhG6vNaouK8EEOp
8lC31jnHGmgFGqhe7PHZ9tlJgLK4zcso/jKqwnTj8csSILyLm1EOZ6voXzimbBmcJZyjgpzRf9/6
IepK1XwGiaz64m1BvnyDKbRLFMR/It4DFgymwYYvXTqssQfeKXdkf+hAygtT2Lxtt2O7H9jZFmD0
XVHta+UGxIRyNP0uRKYEKyskkj6F3F9u6DWkJnipYeFgV9vnG0ep+VhOKaQ9R2WkQXMv9w8RGXpN
1inPfaVwsxkYUF2INxOA78TVs0dcoKDY+q/6PQPOlxwB4kbuqCXyWfwCsbgrTc26PKRteEyPMAAz
qZaPN6oU2We+MFJu/PN23EWSoFaa+cNNqJ3hN4C3p0r754cfIz9dGrg05XnB11xEM36/bX1Q8Dpp
8s3Wl5jkJKrq2Y2Y64IgIAULjiTiGNkzMBm1+nLjU9bk5pVxVBJbiiXnFRuPhnf5mezr9PriZGdi
RByO4ekjiIaLKTkSm5J6MtYPNJcUmnIjp5zrJrASCjSRg3gk5V1rE6elvYeW1OT24XIRwbiKc0xp
O9exZ7leabyn+6cb0HEWZAjoQ6DaH6X1o6EWlc+5ELfXfhKqjeMJ67qpPQ1K8thfvG3/ZxolonJZ
p8cGY8k2FVtGME2DivGCULb/HTyaCcBrBUVRDYen+sBi1kan4ZuK57nbVa/6o/jHWJ8hXMqexA2X
8AbmANvmluK0K8A5ZRWDYcy+01bgXR8+zlcz3HPuTBxAGlt6FAPkctSTGb+tMAXCIbT7xJE9unwJ
riuwvB9cTHMO8b1Eyoa3Aoe+UP1N4ghyx4iC1NqGG/6KF+jVwMB+zRJIg01RpupYmnAjPzIacKOH
615mmUNwoFhwNI4jvghOcB2KYMYbiUJEpeOjyp/XfMd5cVoDPTkEi8LSII73qcKNkx4fLhiYc1ls
3kXr5gmiWfTAg8MvK4BbRvZEHQZ2ZSg23vRv1Ol1pgjj0LUCEO5dfKPNnaRotYmf1WnVmJnPP40O
SRDuaKPDQle6apEmWrya6LYD3yCfOYkccoIlj314YDCAOnRIP2ApkJSiPV4TqbH5JRi18/iqFIaJ
D5O6KsXVpqXSBiWqTviB8wZmXRIUuGUnXKFI8IEGT3MMRUKLwnQnhVuF8dQPAaBQuVS5Wy6MwR+V
ideaUkJtUjOpChHhAgMnZERHSPIodW3+jUss4mJF8CCPzSpkEnYtitSAan2vWaU00YJZdIKOW/WN
uegCguWVr2EaEUAEZaewKUf95IxgQ7Ak4lIeJNOCXwpX4sQk29B9KD9Xm9duDqwN8p3rBrxgBQXk
IAtC3VmwYlICsttmyj3e9lK7u8iaV+Yh0EDttJjQug0euJ6ergaiUeKnGiMcCMRIccn2ELNF70Xn
rmH3/SRAoN3/K1HP+csqfdVIHnocX40zN9cOTAfIuNPbgMwXXchGOusdaVMlpxnfAYOwITOqQc8L
TeeqxrAg2F6A3ynM4+cJ6xA4XsuK1gYSHznMwj3L0KIUDK8izmS7/SpmXcOyi8G178CsEHDInZmT
ZRYZhv5S57F0wMtbjNRGq8SN6RLEe5Sc6ZIm0q5q2EAuoyydUaV2VN0hiIhR1Y1TJJSt5pircll4
1+OieoIk7HW2tIX7NU+ZjFw3UiK4R2cak3qUE3RNE6E6XGXIpoKYjoxGjuJcsCVUDY36JbqnO1tW
sT8eKxWTDmwkz2CltT/FTfCFkZRqU2K+QRznS5RQzIDJRrmFJvuHNtGOX3GtMW8YJD0mym9saKC1
owwH6IfP97DRqpwiQUuvoEkAq+N/Psn5gQuo4vEufPlyRFjrsU9GXcgmnLpLDhag4C0m1bK8jVKF
VD/tGlJMrrUAOj5WgkWsIyNW3neQ5OKWaTNVi8+50q2PP6zbDZBUQWA9jQQai3BXPesJ6UU+wqx/
B9LBe8ag/7mNyYLm5UdxoTWYEr5xwsLnmvHW/zUTAxdip/NpEC8PEBBBJfbqzsiywD9pay0wC2+L
Y/IoMcY274eLVKNYUxV/OMtHfe+B9EfRiSgNeOhL3i93qgfett3mSXN6o6N/8aowf1psVed6U4rR
wmTqDYW3htybZd1uGTTMK4V4sg9rtaC+mLMvzuU3S+NMVGRGea3YT/u9vnrjycC+HJWMLLqiVNju
UYxc91fW7f8FqL9Ukj8EFyd6oMTkfCDcDS+3Li5PhXx9tUik23aF294JGhsnZbWeIm/+SucMKvNg
YegiuMO8OyAvrhzbNAOkZMGLGuq0o12MlcEwazD+UFvqlGSIu2aO+oqVDeniPbewinHUzplUdICt
bGSAqvRRFaz5Zm4UM3iyDtgdAr5q/W4wYNsDQkPS13vBZToBl3/0LSZo57jnYu3CbhvxJPSv3mLw
QkmCUQfz15je+zpC40bUW7YAb2lGmuJeZXuAs5bjqMqjOPcqZdYOCmLFeTg4I6MQkbUD1rHwMcGg
0P4aNUntFu4SO2F7OwnRwJMGFIFDhglxZT9tLv2AOdGMrr/Slp3AdpHRXI3qz/WXpAVO4JEsf70z
GO2af2CMT4BB2mg0jGhlGsspfJmNCYqwLh6NWw+R/o5xRy5lytSMEDnCR0wIKcBta1i3uWz80BeZ
UJZYuL8tlOVUFhVSNBK+FSv9GkiUjeqIfIdzuEl6pCccXRZydNrLVPKrpvU+IlsH32jgV8Hi1vdy
aSZwAdzcnhhQEFZcnZ6YBtieiKkOQu5FYv8Ut3Ee9NmIpUkbRNKz2rbiu69FAuQVSxWzM/rF9u52
22Gkx3QaiynF6lP5+WlwYcnCkRifw+vh4ZU7fxHrjWCqzD5+3enALJI/Up8iqjXWF3rzD3fvAped
5Evu3c7U4tqSbm1SQJwGAhyOQRgtHMTer93cDJjMadRujqEx/5UWD9NeZwFa0aoDbZG/6IGLVog9
LVvofXZ4/34MqRG0jQIBltEDb4VBuVg3LMTqaJ2bFYZwLYBDN//IJBQtcj2Aj1b0Lh/kDrG3ahe5
nuVZlHgX2RQx6cj1QUKOSUwfOSBuLlVMDk6lGEhXyjCIqw4xtPL8IkCf2mfvh1Khs5QafRgiJ7Ss
lMVm2h66zo8KQioMtxG4gQM73YegY2CCddtD7JXjfTCXNP05c4tttUDAD8LLAPdecL+OfTIDAaOL
dgiy5ropwHi97pTtWvQKBrYek+HbO8u7AOG0kOGR66DkxxKDgqdIcJQBK5QwRUSx9yiGmySaYu6p
dS26hmuUBR5fLoSsZWS0LP3jZAg8MRVWWcdohxJvOqT9khuhM97/HBr5T+vyf0g0/h00hJ/sJ4Ao
u5Akg1NGMlrBcDEOmu/6cf6dWx5IJLe/8d+CIDNYQh5xYj3PnEkxASND/H0oPMr9zDWlHAU+JPAk
aeQ66jU5pdNl3IUqXqcgaDiOBflToT6v3qE6Ctj39JL8vVrH8R6WRWR7NqpWqOjLD7sL7e7qi0HO
o9bBkPm10C+mCPEMqvPLIvxnfo/1NDeELs9qSwvP1BdeLZl04iNmjohPFMM7ZzSUYtBcKj8IMhWX
StbntQUE5gqDgXpRsnAVTjKq07VOtVHX0FrqaOk77yV0zVA2x/kctFqc10t3PypqfologboFIkPW
fU+/kpw3kKjabe6rxLmLmzvRSzX14ic2DOCp8kXHZ3fkq1LrnqyfSbVuw3b5ZcCeyOKo2pC8bA5E
kTdoHRTZL3YmIwCbvgqSH0woyLiCUkaf3jmikpUpPUzimPL9cynUSDAvXtnldCkaYxoznIZm2yvW
4Z4iPTZPZmz3j1ic+DrTThfpGyDLr+AwhichqvswTH5Xwfy6bOYlJKiMA4uGE3FVLLx8/X2cIJHr
JntmGwsq007nv0D6BGYQupcs5Xf2mWvj+0ak31xMhN8ExlJ1Se41i9G0MlXvTnKSNpVRjHtBs3fm
e3XOEvovdgwSvXJjBCNAUnSSnHMd4Vc5ZEetP4sdt3t16RWxJMn/KSw0px2jIPcyUxMZYHKqlgf9
MneKU5vQb3yYFP51dAcRAJ7pIPV8GNKDip3s8tYkwB598on8ZZVT3JGblNRtCBG8QEIAtAe/tgeU
3/n3+mnl+zb1+7OFfBvAw1gawH/jcS6gxt2RUXgz/Oai/TZeVq0VdZ4085TFAdaZao3Ax/eVk/3b
F1AW9XM1+Jn4Nsn2738XvEHCwUw1LBdebkliFRpNpNr0RLjXY9Ra2w4GuY0PztYN/4sSiBLAyEOe
NPk78ELgILdaTugbUcqjlzBPKBN5SLNx8AQ+5m4nv9Ns1pSpcL17SGkAmvOT/DTi62+1WmCAbtCx
v402C/BXT3hp0xY5CkIKigUiWEJP4gQIRTm7dYTt6xHKfUAKEBzCaW/lCFBIndc4lV4XjrYCLLS0
5lg6kkLW39jUi+ggM+olu8BUIQjvpWBhwwmalPhAqzZvFad4xyRjiBJJnPBwYdlKXKNKu6j8msrZ
4yY9fHMqH9YVlmR/Z87xWRm1VAzqh0RZBt8vkVptt2XOhJUREB9/9BjE3APEtk5DLNCTTafL30Qw
5z5VcwWx2t+qIR2q764CkJrFAIN6/zt5vmpR6B8Htwna1aYgyYqHlhWKZufFx9HLw67ByX9Gwr8p
I6YYXr3LQjITiBOgZbdxpkYtLsBLF0/YKv6cN9CtroidzvhAlzRWpQ1Hl7QhLi1hxdlSinl5QzvT
kuowxY1uIVfCHP/vDsvFXrRjgzc42nt5Hw4nS3O0YJVuy872PI09wmeZFFH6LX/yrYc3gr0G4Bu7
fIN3gxTAGCumWZqw2EIERQwB2Og8BTtj+bFCA3ROJVw0Evk3cyNySA3qgVSkxyq4lEG4DNklfeR2
XUmMDDy4VCsi8AlVVN97UEF7zt4sJCcTh8Xw8cbxQChaYTTQ9gthKUPJYKlJwoewC6ll8497+n91
f2//izX2i4zjF6nZDU2j0lPX23YDNoLoFQCiqAQ8d7sS2LVJP59ybgKgSZ3gFaQ9380sLrMbu64r
MG7pAWniMWbSGCwtP3aVi2OKpt54xzhZoKx2ZT6eYIgZugQRzbZUg69f5eABye4dNiFYhoMrJTUF
DwQNFMlC2osPpzdtZqYQPCzgh5aWcPW5IhSm7dGD0amIY2IfIyZ4zUb834Y5Kj1+/deZB5zp670T
UwdNPYM5TjCTTumS+dJPm7Pbgkd2GRypjKdXueloxz9xGQmtuj8MdyZgYFQuNz+jMfLma8Yvx4mq
nBkaaa/GGzOJqEqGO/VHNHjqYMWD3JjII5s3He7qUvzw93txs27yzpCLdKALZfxvi4ZIASdL9xbX
XLL+qdMSp+sUfARC6Y7isDPqZJqf1iiNGBWiG7pbecZ0UQoY52jHTMzage1CTB/RDlR3mhN8jHEh
yqWQ3IYhDGN6OMXUswvoJEd7enuMXfU7zx1Q3atZc0phnBQOtXkbfjPMmmrMxzPUY/poxlccx9sJ
lBcQKo4Y5fmJAVbygml6yxu/1YuN4VvPxWGsKIVOy7i1opG5/m3U6CPuNu0gbsUswkhQFLTLVotZ
kRgBIIwW6aHOjrJJhghn5VwebOfM+mWsh7C5hayUivS03V5BJ8YQNqSYTmNJoQcDrmCB8v3Vjeqf
cD6TfMKorXN7IEzJR1f+perUsbQ3mm5YUEvpxuhRiqnhYhZkqCUAVA9ugPfrQNe862DxYCkj/Ne4
bCrrOGH9upGu5ObYD8hETlJ1d/EMWbRTDgfHXyPwP3krlHcdpWea1dgN7T1VYdwR+ZX7Sb7Jvdpw
Z8GC0XaPA6A5h0avEVMzn5d4kq+bJEfE2NQJEghSGLu3VCkPXbweqo9YFvGM3N1/Gvs/IVNIlqK0
7fmVh2W64gpI6I8JXtwZGED9g4w/JDm1OJcfKPEPIO9Ohvp9J2++TS+PQocCqz16LGBPexuzqlN8
+/bZndpSz/utY9CH6s7DVWAQR9hWHZ4XH3E+C9be/wk3ywX0BJh8Nef8plX9MSjy9fY97faABDra
YC5mKqwrpHz/DTtbfCRuPzgXgqODNcZPcZeC1htVq2eRubLSvZMM1zj3XasZq/8ZOTXyus+q2ZX9
//XzANRe8p+fOkdbH5OhU83RQpLiHGlmbtnSyglQmCNPm5XRsKxWq7Xsu9mKFCW5PEtON+qCdwYa
xPB0PyZNVT0OvTsSIrKKG1DL5yFzk52MrxlEMC8Azq/LDMyi3WAvcFZD3qw74/2SOYFLNlyk1j/V
9pMxBArTiQiMP+f+Il1D30k80QDv/JBuX63PulizNXNDYCrQMG9Dj2IjB8zTCiu1MwMVSX57mb1R
9skqLpKgth4sOhaKTBgB6dQCO83Xbe0PBNilwaawrsrw5FwsWV9xoQySljs45s34WlSSJanZDA8M
ZXrp80AjnGUvTIXwKlMDCQS+QwW+xy+mnvSKT3zEY3KuLtQ+v+fffiv4vXzbEGCczf6Y6BzCF1yS
dX1ntgaF1A3BxZdWRQoLBWhBZfXZ0pHu75ytSRvlJCkOQFdJefIrZ8PH4e13LMZPLkhUvC2DH70b
pthpUc6pqOxsBhfepvwslDyS8qv8Ix3u0eV01u+nweJgrd/o78u8fvRbpqkzpg2/3MAB2s7gyXzP
XTDRi2i7wQVvdPd8d+qjwhNknPXAf+AfmMWCx0JD93i+yCZAxUeyWzidXSXHy3OCZBnqcJq+UdaR
sWsOVGK/IgLzzVCnVPM5zyPrnUxxl9r6gfGRiOjpyhc9zj2pbIwijl1g5MKx5K0Bwp5J6NjFtBrQ
6y2NXyetnAlsqV4jFbBKCIcgJP/OM8QuAgrIBSveHsrGJfJlazrd/AWJEcYFeA0JVnBJHO6/pCtr
5QldPDECmUOyqMMJUN14DeVn9nSH4DiaQszdbe3MuKj+PRi/kv+aMMHq0KZp1sxSnT0prHemVn3t
FJh3uS+FC4WRIA2WmFkxLJH32H1zZG8e5PNPnY2smGISyGM2l63bJgGrmhrMUd546RtrVELSGZeL
B7GXFjHgKUE4dF1xSdaVWcOhFTcVyaH1wMNzUHOMjLPpkPD/78FfKFZ/HjbOL/5qqYeOG6u2bvTd
LjH3AjiVC4cNdXeMYH6tySb1aZg/yDGffxv/b+HKFBXbdiGEx675Nl2wRMjMEGRrqG+CKLb/eXDY
IX6JayNmbLvD5+mOeQHhciBHktKeZabEVC+XlnaZYWAtO91hPiDgZFTFtEAG51TeUaXApf05uc8Z
s3WqtzqhuArYxxX9Ta6J0xxy6lIvDtIpF54xpArupRnqjW4gEd+NDh5Rx+za+HhEHGTtw/lV5kND
eilEhtQGWH4WZQYJqE55zK9H4WZV6IYOowKUgQrzCWKV2PzErVTIe+YmqWNjJENny0Nl8sMNJ0Ya
F6iLdhQkzaPudTi1JkMPecdqD6LpkyKueCUyB2IlTauTGOnUMq2jKjDDlTlrr1gwMZ5dgWcLMHVL
iMRSXF+tuRVbt2CaKL+eKX5fcUe+/zkmbFA3NasPxtQzIzriSp3A8hnTJQ0UmvEBRESZwqvFnrf6
Wm+DhX08LEm2YbCmLCO9/3Si4U7jUhpVGVYw1k+WZw4ERsSMfJlqHGQIp3tXTr1Nt5fdgRrXZBa4
WviFa2tXlzi6OUo97HSdWKQBlE2jEyBRt0JblWy9ZOiG5R1i5oJQ5s/yxv9vyZx/KTWsDbDgqRGd
m605ai7T4pBJ4gIBu2X8+iaJkS+gTjtdCgE159AppNmlG23Uih0+x+b2E8RTSlCYHucwOCN7+Kdk
9IwqGd/GzsMiR1WCGHady5iY8kTcYb0+b7OYebELwF1zrAqAr4CqMybff6flT7q2UT2oFk1BMzeT
9vLBmarmQAp51SC9npgBhsu2/1NgvCQ+m/Or7ZVGJ+vItuNIvH79LxoZ/9Soi3JobqQ4mZy+E8xv
QddissluhHWiEt4ipmIWb7xzT03qYId5uGtJchIawhPSYcEvS/XA9lofcB535lTfMzLesP44j8EW
o+Uzur7+6Gvz6iFoMzQ2sOikhwY4XsdV1eHXZ86RCD7FfQ+tH044Map5ZSzebvbiy47atkubV601
+tH/ZI7dYbFCOBHufZnsdl4Mm+rFsl3vU/Uyd71QJVnqIkL2fshMCdMRhBiMHx10Kv9BTwOC4BST
l8vC7blbDt+ae85C82P40NuT0g+5zzzATG4CiV/eSba0zAZ9VAhKJ9zzoxEN+w2RdTXFjWjm8HnR
pUb+r0c7VpahjDrVbckVsV/zm5EF3nNw1bp6yOVI+qihPyu0lJ63EVjB1w9mbPmsyMDyuTsUSmR0
Y6VIwxEqxYpA6Bp3uHXjY79XxUBQ1zisV/OfrrukcRyJLqmROM/MAI1T6Y9OVqNsmQvImsAR4M4v
X3dRYwnejCSoWI7LeaU8LClpQC9DqbByx1cFYEE16osGmvSc+xN6ecPtBM9FiXMfSRgr7/4W+LsT
0W4VMZ4hhW0BljH4tIPZnhXkcL2uiKPFk55qrXTEgN/swN2sW/Alg4THKCBzR8JidcXRvPgNKlWz
9Fa6or0CoHTpHyWnY22PiXJSpDKTp+sTzHYN0LJPwr8PklSOLagAQnof8YlidvbYOkfQjXzaqDc1
wlKdqpN98CmufyCzfNvpuP5eQX1O623LinhkdhDV51A2Ges8CCw8hAKN4trEVdXyILhbY5+JGINi
rerg+GKh01PaP6i7UmARgbKzpOeHMdBEUCc1rYIT5ZBSpY7dbnwYjx5l7ask0mp7IMfZKO/UYDmC
eNVzwSI1MtXuD9j3TiyYbCNnm8Zz9a+GI1zdkWmZ7uO5Ir9H/U5X8MSig/UwFpTn+YP/00d9pIST
4A8b5jTb8mB49qhEGXa/5DJ5Nyzekf8/gV5Ytuwg25Xcrcg7eWnglyGMigEU1qV+FUAJROy6uyTr
w7kAGp4hNEoXnvXos/bVnIvfBcDgcMf3ZKmHvdgGhTVOJlfpbo92YqlWPkrvTVhCtIotRS2uS7IS
JtUZoHMTgxNZLziGc/5oPvlYqxkrtZPGSrV7yV1d1ncRgKrrsllLE/b7jv92xGXAg4uqgAMgXcyO
OBcGnlw2FgwbFv9GEhI8TP3SDIXQf29q5W5JdU512Z4kDhFBesWCdlx9U/Qs9r4S5gTeHBlQ9pjZ
QgLSZY4Bk+hrfc+LjZXHk+lKYAStv4N8O3CPMogKbVisOkvwAlBlrHNP9wPnIh+piyw0ySY/Mw0X
xSQ+rjqOqKSBCIr/8FKbFiz3hftoCCVRzbKIuKOgmqWwlxK9qPmgqluXxhUPa6vLyxHQd3lMYmVV
Z4woicYgrbAag/5RLEpSirgxehy6XBt4BEqmc68OE1GNdl8H3/C82iskcgRbNBorwokp6nU5MGc0
pGjnERXTpk8Dxr4yWTt5dsEcYBi9QWiZ9uwkNvUTJMEm5ObDao3JdaBpcOn3ooxhRofM5ZBvlgJz
35flLozHjmTdUzAl0BWgcXdOshJtJehZcUj3ExkwuWjjrZ5hPHgp1bJ1G/LpAcecT1KnhbE6AXa2
cgVB0t3Ecp7pFxdsLHJYRKtc2s8yCPb10BuLf7F+Rx4acD/Kx/lbtETuic76hz3fE4gOESQYjvRf
+ZWfsFunut2m22ncUOwS27x0wLMpbzi+zkPvqZPvS9V1Ols2wqZkl0pDuPFyhz88/8s2RXMLQ+v/
9utaNlkzBa2sUwbe2xZiUxhsJHYZgXFsl2Kxg87NzEbGy1wD9W8JTF7Ae8IhjMonga94kxJO87B8
vUtNJNlLKzCQqH4COsYG2LoDr7geTXL+MfH6r5we1cES8aohOj/idXjw971MplrIOF4wdC/WnQUD
mQ3GZxXmhhEvY588UFMJ5C3lREYUpBRVZolrD9rvQayEN+lyTtCyF9FNu42E42sHzghV6FgFj+BZ
aO7FGN6tvNJ2n7KLPQyOOTMg7qG3SGW6Ym6XyvOkJF9dtoDLAUnNA8emC/BMa8JHbY0DqrOGFmgE
zT8jUSblFfT+64oSaFALMJpvVvKMMNShBYEK4Y/iX0u45POuNBUzu52qkUMbl3sWbm7XX6aFLVta
FNacjHVGZuBo4/++8TR+hEQavsaRX5+xqDr+0qmwMM9XckwwJamv1fLL9DHVTxGDgJnQGaAvGoi0
pD5aVI250CmxxkSGqcVGzftISfxI8SzBr6dB0/0z7x02ntK1glm0lfiDcB5jBec/GmnStqWKZ+op
OjN6tb7RbZ8+0NEEsP4XE9QabqSK/Sz2EYvibEVFOGzRM16BfkV86TbKqSy5FBpBBKN/NVp4n0ri
Am1yqEXoe9G2Wk4DEMvXUmIOS2/VDggPK8f2HDJ/nVg/33bHKU02BJMVSwitqedSl5/BKl7Gpt30
rxGyhmRKG9+OPv3y7TZJbqkm7LlV2Sd7Ix3x6UlzsG82nqPmYfcfiFxc/p8cjKuinnRUgOsdIlr1
x7OjCocKEXOIx0ahEbbkAu+qzxaLWqRQvbr9XbD5bUPyFcytNOulfvFDcapf8/RayqM0vmhTIpbY
D4dWlpfeserd3xKQqyCeg6xNTXWrlYCo2ZGaMpq9Y0Al/fPiC06v5zDhPryEPo2ACwMLssV1rI//
xYnz+0vKBo6YujGERqaPkBaKPyZzABa7tkhOA4FxTulgW5oOjXmG9nCzVXRG6zbJ3dS9nfNrkxI8
PfB/XRZY/t2PVwa9pi2VRWcisgk42pPXbnI2VqWpF7NNy//yBfoYlMK9iE4tJKhxrvAcpP19P5W3
hG0hOl3pyaOVVtir9UyFmOnYJePs0qfh0rqZqaSltkFjE+SYyDHzXJdrfugZNcL+HjevR5Hsu6Y8
MsHrwkscUKW/OHy0G9Qj8tTLbzTTiANXG3kZjm2/KzsIBbOQo1a580jcfZz0OeO7CyN3Cydm8cNR
wM5q/5/adSrRXRrvZIVXTZE0T1lsI9qAkNNDImMmLxNn5iG2f6GayHVRVlputQUt20DjR1wlnfxk
ycEjQEwuzQWkp4ce85LLj1f2XWFOO5mGWcc726Ozt23xS/hVAN9+acLs9/HuFdAdb/URtwbukrb9
XWKRGGul7HBGBf789fsNdKMNoqcYlXO4WrpkGDsICsThmE/h65okFhAvJD4K0ov4N4tSqRE1RItf
SAlEnu04FwrTCgkQfvtwABMVL+jSBDUhsD80AhGRaXevUbbqDu2s71fE73X32iqIPmfozuIxFBfV
hPtO06xKCO1+O2/tABE5WJ+Z3SqKD2BjFkXjHqN0f9nYrVPgEcwfEsI72ErSsX3wrgTWj9jD29OK
TCDMm4DOfXubrF24AnFGjAckxUohxRLio83CuawMIuZiqCHUOSLzisZ1LHtL6EJ9zxfum1+cH+eW
nvAGBxPnWU1Rku+gnyRDSypz8I7BXHW5SkihH+wsIo/LVqsRfkyvV0oU4K7I+SyYqZ64v2mWUQYt
CuLydm93iZiBN4d0AF5FsV//xfwvlDnV2BxeSYF+/Hy/FLzfycL08ht8MLpSCXph/1XlUjwp3Mkv
pznAAyixJcgPZlG9iXLPwdCZ6BHIWWXSPMhCNW43uK+UPBin5RkPOhkTddJKtbOmeDqQWH9bzD1Z
dm50TgAUgkklPbceYLpPK4XHRFqNZuSd+wegX7HXrNxVgPUtXPmWqox1hRxxX2vucJdMs5uU8MyB
r8JHsIPjtUJnVKGCUEUgFbYxbdGqQWAp+2PxUlcQpvFXyb519FzAwlzIgn93+S7KclcDImGpxAX+
q5KgEXJ9v7N0jieB/Pp2i1J3OIYXkERLcPPm4rfzqJRpuKPSLGSAo9NA/U98ME8Sz5UhtFsA+/VF
u2Tq68Q7DAwrjvvgaKTzvLTAxxPfSZYo643IQawuswucpJId80fIICOIARnvPqwl3vSiTuKKP+6W
DJRImsw5E+rl2ZPoMt8Z9b68HNVXZWDzzNDOrGPUOAlSSANmWsE+yzZslfdpgQGREWZFlHjAZAGy
O4m0SHF3CWrFuqjfdqxTUSqmI1ItqktvN83v/6kMRJzDFl2h6/TfmPNn6/x0ptCnD8yAunaK7x90
g5fU1JDlf9BMg5SVdaUJB8F6C2UI1zMdUNycA+anwXI/KK2od1T7bvyiyykqjoromYBwmRHAF2IP
kQ99ZZEFO2omHtRetivyFE/vgWEwxM8rTS8i5m8Ch/tnyEMI1+HnXfTI94vkQGV90HXJAzfzp3m5
xJUw7UhVUJgdo0deUPs2LYefWhuNYExqBBEVSHQ9GFmXT56j1WRfUXLgd4QaKgiprTZKDJJD5RjR
EU0cP1E2iKhQaObnW/yKQSVA6mU+GKqcTND5Mbya6ZGFXZMgUFt7u0ANafaTM8DNu8FpkLfbhn4f
z6EdgxopNEXQxh4hR74uoAWtmh1is7/gfgG1lVUZ3p63V4Dmt4YAfIVpC6X6eNlU44dOGTHKEeAA
b0Cf11KZdceEBthc1esrFLQQywQZOGsD0LD6+MyShqY4rQsisx7L4KmmfGx8c19kvWwd0oaLWXMC
752luKUJguQdf8S3ftmSEWKSY51LjN4dY92ndX8X+T6R9zS1PjniKVAvFfFl05lP2ktvHbf7Ckzr
ra0YtMa4YZwYcyfZ4nL0+bKpVjzXucbPJJnVTdDL34taL6+1u1yMTEW6HlY5ApxCGbcpbh11hOxy
Sjzmt34TwV2N43cntupGeawYJ89XAzPSfjiOkJh/c7MgzgAlO4rrgbjyL+kielE5eIbQpIYHR8tS
w35j132WxY+1j8//Vz3KBjSIkVr1ftHpe5XPmnyZQV0cfjQvcydidAgCBuJ0IRO7bTSW05iG7+Ud
BrkRsCGwR/LUJZ+TG5HE+cEt6u6iAz8+vSkcWeIKxTAYo7uxu1+UvjYF86uuKnDkN3dauBe95r97
wNicmcILjksNDZ7VvVQIR/nBqFSdD6JBVt6L2f6qweW02uPb4Uf8Dm/4Oc5HP4PY6vWnYisQ4p2K
qa0YOkpNzYGi8uFjVl6J1y/U+w+M0qfcJflKqfKIc2nhSss4Jc9XsqhIyAshr3ScWfoJpD0YYAly
ETXeN7XzdwW+Vra4IKBufb96BvTSDXPWFAYpPK5UpRmLdwuDbzanlhIWsxoqyhEZLfR6KLCKQsGS
BH61qevJlTjkaoyQueca+MHSvfiYnCZ+D6UDvBoA0siDfejjtoJeKLdaXy3FrRfPDlMqL6FwXHbD
KrLxGcoK0ZH0Y/A67K4VzJaXk/zwPDGIS4TWMWwGcMEUkeuqSxPQDdNVdjTm7L428N38RdbSH/+1
40nSRnocVbninxtnmyuV2pEAeXoN5A347rIrqPe8WcQ+YLrQtMUnL6t9vrZSVdLTUi8+ZTvzpDuE
168A403yam0pK/g7q/gQ80JtOEIfYJ7OwXVaecnKx1dKKeNF3/p+k4WXQYqOHQ9ugaAI4PnG6KMH
ID9noDO3Dz3OiH2w7IjoZzPqAK46TDnuvwm/XvNbV7wUltOU34RVOlU8yk+S4o0QopIdByWZvO8F
1BuTTHpWnwefQ5y9INqteitg/wyYsa6Y5lXU0JTAgqW6MwxrqZFxWTUsEw2YKvr0qwicxb8idKdd
i96P33Q8eBFqx2fWmwuTCWIycTLQF2hASWP6HTV6AxvczZ0gVBO1OaOTeMseHPnGa3OfayDypH7s
86wtTZN7Q0zAkmMI3vbDPA73eNZHeOnBJhY7KoqcaFP8MWS69+hIWtZeT47PGt+02IFdbPLC7Idx
XIG+1gaklqGy29h858yq6tf41BQZgrL20Of5NPsnPq7htjHTojW3LuWvSuLXpdF/YN1T+bdcbpnk
ZfftZ12NrZay5Lhr+Cppg38b50Z9SFvZLewV6u5MAfFV60UpyRjeFpO1V/dvZjtsGnXViZCh/3Xp
FxEfsAHFyXEYUuei57/08HRb1rAQ+GfpfwEyFBsG0tLXRwuuaaskC2h0BJ/Fsh6G2nNbbg35k0TK
dbS3SfGhFnZJuyKMe+1NVKuR1UIt6q3qyJybCbth84BiiRN0Ak3Ji5RzKLhxAGDAU0p9OHqUk8cv
ccOp4eP/5yxp4vcxjheQ/bR3nvEsed4jdROkvxBHxQtF+shfpvf1udNhb4/LZiayIKgjs1/W8QaX
X14BTsjxsD+9WCDzPBOtuEMCtnSFnCJiI2cl9gfO2OQ+iUguESnneKsPDkNoxnUhQqns+Si9Gi/i
OYrisj5NXit3aJlkv+W8lmMewlejkxX1X/6spzXRV3Fv5vXvdmSsPCQBWKRL4YU0H5etMjlzZ56Y
B5nnpqvvG2kRllv03AQJGhqPJwYvc2z9iVc+S+PF33r7xswNK+0CjAIH8FUplruSqNecCF0mrxt2
Sa0WXwSVaGBQF5Aryvke05s13rFzPRyITp/a/8FEF62NZaN81/1vhewYDNOZhbYHFzgYT5h7xmAO
YD4elFEm8xS5b1ya0SEK6/yAzKp6/mfaZAaqpzARwVXKZXllcYBjhOWGvmwasKscqY1Sq3L8ruHg
C02ftfMyujb/trnz/gPPMjHwQRdgCLQcKiCviz12JYBg+96LnLUKwF7KMKW4jiES3ppXlYSwRcu/
M581WE+hFo1Bhq6nSu4j/BR/l5mUvkKwwIq2TG+TxDxwIGypi+mxiTBeeIT2o88bWcR1PxjxJwFv
uWAvC7TJyItqL2lyGdM0rzPj5ElLo9xneQdJPZGCr4ijSW/BnddLXUcQIldTRk8qBRm3ZR5dt5dg
hy9MeDm4X92AVmyv2RE9RUJNPb0DZQAxW3b6R4QcTr4Fm7RI5o4kCLqUCjrDg+FKQi/SyVXvJzd5
iL2JMZ0dIZaDC8dQJoQSQ+O2vaG2VifW7tVFF/EUM8oIVDNDx3MdzqdE3WS9W7VBmj66hAz7M6f4
ssYCoHezCCYG3Ms6bdVlBot7H7ECwSPbA+QWK1E6L34tTxH2UihjCz2lA2TuZsE71aDHoe2uz+Bd
KhvylkwXc2BvSBgcpDaPTnFA1cy9WKTmi/ip73jBe7iqT4eKyqGke6Z4hwZQGyNN9COCdj34Iw53
xXkukyZIImJw/jBUWGYIJEipiG2JXAFftUhyLIhO2uiG1vfaR4Hl9tDs0Tp3ZpFBfT3oEqvxfFwh
owruCCvtphcGNIGNZeWSKtEDJ8o7cG8rmEUyX/Eo4fOsMAna77RmRvWsLH+gQ18KSRwKfqrlcWMw
xkRu84if6Egc4CtZAmtdWt/w+D0+DBk4WWTXMTk7/mVJ2eccTBLb1AUjiABgevZxzJs+jgLZHDIH
hb8BZX3QAIrceW4lRw92sh/20jh3A77w32/nF9Scgi+V+CGiH7Asf68oraMBwFEzYxicEYTsShwP
jPpWnToBxha5QzAW905b2MoLX5t9Pi2eNRjVJWXZiTeQa4h0osX5fefStxvQxABTFvZRAY2GwO9e
kfF4XS676d17TrImkICP+uKq0dnR27uis4QkyAeRjVtTPbAhRghdhbjoO1hft5ffCD30bp0QtEqn
Ja12yXnDHB0X4zu5I5dVlnu50Lt4QRpr1drG1PIOnj+y3nGBMimASEN5b0Ys/CpEBn1p35xWTRbt
ZRIFGry4qGgvza/3tPHQmDGzQ2924+vyRcCa8eCgnDsrqdoDlLxwFKl+E2hEu2APiUYyckCFpKki
+5MZdkX+39Cco71ZhQCWGmKrYgfpDDpDDrE8WrnVQZGO8n/wx3HEhkK1LmOIWh01s5byJCzCTlNP
tiLluvSPpB+1Okx/1vpJRD/7AbdduFK7C5kVALEY0uqgKLq25FmZ6Pd/S9Ji0WKrGHKb4wxfsU5O
5nyPn7/kkUo1dguB9ipWBgSMHGhSptaI3Sk54Y0XVVWA6rrjhVQkSiNDZ6h23K0zuPPWePqWpPng
ixT+1eRwzbNaulpbUgaleJgEfsSSXiubSQGmdWTlEhHaxHZabSFZEN7pcpAQ7QpbxrFHPxMsJBJU
GLa78QjQRWsK/F09B6UEwtotuhQTMOOa5ObNlV37Ghe4tV7ivWErUky4IQ0YHsfYj1KdPJwJmXMu
rJvgelm7hvHJnWh5QAjovBpa40wSdL4fUkTn52DaTXZZ+gC+7peqDWrJ7fCVihPuNTLFIHiUlzkl
kaDK/Jju18hqJr6Mgy7mFmM4xJO92rhdG/KnpBuCLmNBYY82Lxwp59GmxXS/WSPLWkJGB6hJ/9OU
fzzjJ7UQ32mYb0Yg04BmCXUdTXflmc8HVhMQggGdWM5CAbmdf4HpRD5HTBUb34HFmS11vQyKIVIE
T8GUiACgdRG4oYYqUsoPMKe4WQtpp48j50UU78O/uyRBHrzK6ezdmjtPkJifaNqd1cYI5GZ49Bfc
6KxtqeKrFQQWv7F/c/1cpJZUTCiqbVvsUaNwN29UxVTk3G16Ida1LsteWeL83yM8HzOoPUkOhh/Q
Exl/gZeSyje5p8PMw+zyHgyD+djlnR/mE2B/mkcXj48uIUCMCDKgQ9klwfYcOYdkiVYc5ZASEjN7
/DDoN7tbp+op7MRgmFJaf1ImLSJPeN3+ZRAtiAKUOB9i2ZZF2+Ig5j3j/EdYsI9bLA81wUmrn21e
x0tu+mLu912CjYrRGuPwxanmxtywN8E9OUkwwvbkkbtRtzfq2XNgD/D6WJWTEyPpIbk7yTtWiKaT
mc7uMDsCnAORR4uxOt1wvLq0eDPc77BrXr7A0AkZc8wxkYjzY1Jf468Q9ECZL8F1NbMzHGu3Wvc5
X5ztNxpmcngodZ0kWw5hvWjyXrNrQPT4SJYTc0nU2cFyS+7+5vAxBTWcL64in7zAd+VGi53zPnSj
ax3l43d+aN5W8IOXzRwJtb3ZQBH5BEcsR7MmG/UYfdAk7MauWdUgVQbs2CEoAe8NnWz020NldYFN
RyO7LQBzy5sclY2Hfl8BwsXFSZZqrnaWnhKFxJzwepo2ry8Wkh+x5NfuMQKhob3DYM5cljbXdOU8
Gl5lfFM7W14OF46dGc7ghasqOwS07raJl1E7Mqf31UPTsAjMIEeRFrHMM8LMfsvN3oNmLRnmJcSe
LQJ+68a66XfPFHsk4DdDn5F0XVNi2HN2HlQqz6l/73emSBk2HsN2ey7nTMZ+7VPYrC8YwnWZcJrg
28wTHB70fQHX6xkKyU3Jfiv1xyrDPdwetNHvfEps5ZEbsnwNR7zVQOFK40mGKbs1sIj37VKG5gTS
vL4kPqITV84VMJv6bbGN0JbR8uF6CdPGmbH6H+WOENnqMc91pl6X0kWH7PvlC3AFdVAqFp+h6GxO
JBrkwpjAkA8cOhMpwDT7SDS+ddi/Q6TbUEGULExQ7XIP4ksMZ4HHytF+yb5Wtjr2/PxAkyF1r2cP
19d4oBJE5lp6z+0/SDYB29fkVgkd8I2c//l0TrNkDjXBqDFUXtsxAB0cssc9LRLcS6uZ+GqI3uUc
GzEBam7RWuoDTNyN0UcyOmbfKJB45TjZ6sFPrt0gHlde19ncIAdHyMkV2tUrBCDz360gzlmtHHMO
IMPY/HUqGh2GYbQWz4JD1gJVaiW4uyjXt+neL8japCNR40RSZVHsTCThZgIw96hvuovyUS7fBTvH
KnGc3exTFZPTp3Aw5g3oT0J4pJHVKdZE+3DT7XkgO66CT7qFUvPyoCO3YSTjHGuE+H20UMwCrm8e
Q6o8r5+sx3pItBRe0UWyXi6wMm2nP9Xh+0C7tew8bHOsIww33aG+7yZ8cMmiOA1szN5X8sycRAWY
BEiOSwSrYHT40QYTlUB7jY+dEM2rEbaozJ5ZjKif79EP7zRD9LawGFo6cbQRxvCAuJCxHTQiG4bp
QXkB3maluUvyZlOktfKqBMOlc0fY3qKUF/wyxtTp+LKfgHc/7fvar8/8NAR+fQTw6PcTbQJZbree
Su/Fwlq7CZJnQCWRCWmAdhdAfcV5nZkQWJJpr5M4jIOLsnHnoohu+SLFOgX0PWrZE+Sv0smXWB0g
fr5bsP9qm64VRRAVJnagtFObDlw7/gEXya08AR2qfgX8XCWkiCxl4EqktsGMe5oV3ac73IazVLD7
UUMo2PQcDVjl87j4ArFuNUZxD2HEBhHFlL1FPMe+mLW3d76Ilb9fKZo25OS/OBXMnFktIUFbsyn3
VtUQFSRc3sztvW0B1HFt8h/9X3j27YWJAdSuo/etyU5W0yl/gtr6jZnm/76g6DKAVhvIOmmq12zq
PSxE/Y/3+xs321J0UTqfDal11L8LCdWrwUCXO/u+jdK98zcPK/GAQiJ0ABZx7GMjXy1qZU0aznX7
bMCSNaswX/F1cb+b5qT4MXKG0PBE3REgREmG8sJT6eED7ed1YOqXJBiAxi+y45oGejB9t3aCexF/
EfF8HdlE/Mj59udIehJDduszJkc12Rf9nUMbFVjMFFYATNnm4TOgkzrFdWPQuI0tPXvb6QpNBsqL
cRtHQmyaDemTnjVuUpNjF/ODZtQX0HdfdPbWsSiafhh2Ta6Pi9Xttw4Mdq4fgwrexhMnDUvM4Khg
tiw2L/gURBi+WUX+1usBSB/aEnoWUMDpO+vr40rGyF0yp8Z/mlBCT/ju11BJLiHkpJYY8ErcVa96
6J8DJ0qYnzlvcMCIvAK/6irO6TGfL1kH9j7jeq+Ilpm7NpDcrIlkTKTPesZyjCbCNTVC3LJFWIVb
JRr2A/Cff0Vpfa6M/TGpEWcMoPJ/MEh99zgNcpqiqXZxvWcZfyfyz4nUDdj7Cr7V4+zANhYNnv+8
rw3HywAn/MA78PzpRTIigfELKTD4idLSq3AY/E2DXjfPXJb8SWpdTZHoNKQ5fZoOCpNHBj15H/gI
Xyl3zr5EgYnEqNbgCPx0w2WP0Jp1IdH175aOG7f6VfpCv4pcDAF/WKCRkbuqxXWXa4JI39gO/2Aw
6tbMsA3I0Lqv1ryp26zDdn8fvDgbTqia32z5HjLWNOOi0n8ahXNCUGgL5p8aFJnekyGt4rATbDln
Cil1qtO/XLYgRfekNtpjwLuDfCOfq8H/lfTPatgs4o5GjiVw3hEGjCoEQi7GbbT7nMjhMLWOb+7c
W2QtDLoSLtJHBhWsiIYHOuO6z12aAX3+5viERBUhw2UGlvx8NXM/dTTsaaRgu4Qgp4AE4zcyfB87
ixMyB0awHzQSXYqh8mhuIaqZe/uOnJT+jdzkQ4VMHFZNs2e9C7YlDWZr7NcMH/MqSbxdvh4bkLdL
YBvbITtX7l8IUoZLdWk0yJe7okuv46/mKh5Vgdmfztiudzoy7agH2FVcUiaAbzzGaODnTOqGyphA
fRX3602NRehlHymiQ8s+ya0SL1E1SVkyk09JujHc11FRZT17uVCg1XkMOwdHzXfOuf0UqxMJc8wu
zXpBYKjHY+oJ0V5n2mtsDzhXc+DUmelF1AYRkaRg+4Zm5Yh38DT1cYz6TyZ+8+UL2F22Sy1MfsOl
FOCOmCVsX4nhXzkYD4fqPEfK7SWzpUpt5/DtFXOKZOeCDtNWDLDj69NRYZHDKeBwO6kNycwk3T3b
bn3D5fWv3cdDThBA/h/4NPPeWMl+Qx0+baOykZelQoD3YzQg7nV0M9JkPGC2+iHDfx9am8d2gD0F
J5Z4WyR+d7yXPhNMHwD7i38SrTLaw1HOyseVCouMp5MulTsd6AdaZNh+yHP62jlGl34RMXIROsDF
2Cgw24myP5IzxabZDHdLQiDA90TnEIlnFTcuy2hSeEdKSTvb1iznPLYsTFtoHhstzY7wmzaPA9cE
o/KT3du4nNIppdRdohDrFgkwIqbWfvZhCBL9iGD+M5nXnPEj35sHYOgy6BA0FyI1cdO1cZxvi+6Y
4dMuIHRgIMzQ6tDXCgLZ9tKA2lW9fNjJFoEa5zQml9I+DLF+XDpBzRLd/h2WWeritfm9GxrG10xL
k9zBfA1woSdFMM29DAW00E091UYtKYIHY+eliklIPk6mg7oWsAZLjvtHllt5KzsxiicQGiONaJ+I
ASRdcUpnhx11IVKBZUndJ3vYCmo7hoWp+Xnt0fYYNFuhOX1ySHMVhHhqJIeSKgj1kQzZCSZ3R1Fg
RnUiUeqajF5xlp2aMbg4kFbxlmBbMUZ4oIGqsCMxq9fNYcFEWeQwBN3tGJBmJf5r9e/gaGy1wwM/
7l0TLGB10+926T1pKGwLL8AEVLBGJpogQ/ZiXPpshn5Bg/YynEkLR+np+D1CVVNxx1M+iktIatWy
XVqZrb2OnfH/1i0fnNGwAjkvdNqxGfoRAmhUk+vUdurlaGZgyv1F5GvAhV15CaZuEt2P6DWNH4Bm
G/vFb79nc7P46yCMLp2KvAOa+RFvsIR52qqmaZRKsxTkV6xmj8KAbbdK3n7fxvwXIvQnBpjNqQ2V
z2d1IkcoBdxr64LXNEmuG2VcXwvNSfdrRxwuVQKxaZvIFKbjkEO5oFrnyTdFejqq8cxliMnZMYVS
6M3SRdfnAGK2t6u8c2gWnLV0UkPlBGlB41Dv7zmZ2QZ83TJwMQxhknj3ebjPNqbLcaKlJMm4z7fj
gVoetX2Sb1seoKhBM0M7Ubs4Bc+2EYUXK6Xnp2tzbLulCTxZ0SKaQvcCbKUgiRbNu1EXjDNaWoTg
1WaK8WkJdQeoUGCQqMc3iW6/BjCE8f0AJ4YvS0DkZFacyJz91G0vLLKHTUO9Rk1ER9lTEyLjwMaI
9EfbMBKKbONwMvE0qMbURj9v/IQlGFJAA4qma+bK5bh8uwamroysavV3EaO9yrpyGYgD4UZEdIrt
XJopRroVlYEnVR5AFacPQxS3xmDjFn//v5eLvIhxjdCEzYH9PVmym496m+1iEfo/KxS+ilAdsW5q
hIpO25I2JZUhkD9De8Gn0RThORwpXSBafR7qJEq2vRmd7eNiChhsP1s/LYovROvxAXh41vRcKPrg
vkUMaXBoEVRPZcmt1uf0+7GdToNAJ5g5sTvKX2mnQshOPSiP07758N5rsMViG8CMWOwONh8wB3At
O8Z0ai+Xj/rdAS/+mqN8dvbwNNgxFTMULD3pK6eelsv8YCcg1MG0FqdDy36TOs2bXusg07zQO658
S/4n5koSUSCpmg3Asy9QcrUdNAOb3M6e1I7hWRNrnVB/VGj7aDuV6PiqSVRCoT3T888aq6wq56fM
AkBWGzGBQ5VH6yHlozbWbDN/COpv7r5ZENNmWbIb/PFRf18tQGEh+I+vCo8fgSJoG0OVHMN0WtYO
4l37OYubLxYBoDyHBUBQ7bHB1GnGhES0PYzuI5L7wqBXlwLckPKwrPKICX/VNTrFZ/QkhiaI/bNH
+PAunfk5gxpgAuukhQinfXEtbsjKw8XoYLuXc9lEaK73woRVdH63X1QRNuNp8pD2zlMj65JZ5eSb
f6xf0MB02Vt/K4MDuWvGfmaezX3E42zq585IOfQlxk7CT2afiaPZKEWPE/R3FJ8VeX+pbHHtwmbm
1xvRVzH/LAFw126muD+2+KZPNCbYMcH/hSVd33wf2B3Vvjrb7KHruf0J5j2HzK4d13P6aKH6tLdR
xu7iLYKwg0SjUVxNhhLkXKqwNlif6iWdl7JPeWnriAg5B9XOwksdeiLLjELk9hgcpvxNH4pt3Kpc
x5h7D/t57Oy+lYW1QTcRfzA8SGpLgoroZdiEFjBCjw6IQQJLZHh2E+ylSvl6Itt8S2tIoL+jCZxS
quEytCCtlKq2inDe4r7/seXrru2v9g94gNkpIQOa38BisggkDivpx1LHUdqNiMmQhZRY7W4sYgOg
MmH3nzmyWQ+UXT5P5iYSMLq+b3EeW8ZeQmjItiVuYfsSnxlwyEvmeWEn+9hBXGDwg1M5pJ/yu4Fx
Yi0jh4QUk8iFYNytZWEcR9rrLA4aQONwvLK4e8eJQkq2oA1pf9iDvSWf2i7p77oQFOTy0zHK4q33
sRNypkClDPBJ6J5GmBExRIhn/jr3a564NPRdXnnvMmycD+kUJB/fGZAo1++xCsjT1vid6Kioey3U
jKzCBiUp4YzgNC9yTslGIPRD9MqxkWyKOAQE8UYNRwgheXum724oX4TtfdXg0/MmLOH6D4EK8HNb
6W3f60iUw9xiU/6Ef2SrUpUtydeAdYO3SKJtnIM7lZeH4u2quCAGkMBTSNYN0HEs8qJ2rgKwyblG
GLtrtI4vaeukzhCoV73+Og3/Ur6d1lUlz315t3/iiI2YE/zaKaIhEjYcvJUvuG6gnasc3TWYNYKh
E8f8yk6hEtfih9aaPAt87r7kn6v4Gr75ERMzmvuYRD76AFre/rqDAJPuZOZq+ZIeFE2cM6wXL0PT
3rfWGf/C/PwBqgtYINy9qSSDQLlQEN2YxLPIhTayqbjoNhQ62mOsdGJY9POrN6XavPB6FTBHWg0g
1kOWsi2v/tou0GDak2npEOCKoYt8oqyUn12E4xQJvN4h/tsjA9EmkOZRbxINADJdj4WANEMzZGFJ
BWfNrLMf7D95mRli436/Ehvjsyqh4ho+ndQHz0WOams+rVkO8vyfhXyh72kOXCRyaIK/n1F3N18b
8mGw/+ISRqaDHMp5lzcCR8Mp44krSr5JqoPFktwKEl5ogYGUmL4++NBrv6iLGXxwE4BkPuX2j8c+
a/gCMrMHvgjZIbM7xWS0CUL3Dh2Tf5uDxmt7MpH4+sui6ywdaXB6cY5fencFOm2mtM+K3D3/CbDg
Bj0qPu+vHkJPvefGb5liWujiZqGUv5gWVGTZQludhsjefbaQJPPZi0zTlRuAoRNvI44iz5SE45If
ID+lLIaYjT1BJglSK2c8gYOYcujESelzp2bwflSdg2Nth8qdaYLtkiLFvqPcBGAk+viLgrB6ai82
vT9SoQhHsrr088IvfuHp5jG4jJK6WIynyAERdB70fK5+w+9xZTRMbNd0A44zsjEgWLqEHE1BGbDy
lhiBfsf/FntghiC35jsBv9kPaAEVkpkAAtEpGvRrbcJvdVYom8OCi/7cUs9hWjwbffGtbjMdioP6
EETCEHfuT84Ot8ndkycfw7TqsyD9Vg56STnVJ7/Gs1oxXf8usoBKM6dzJ47ybNjCSgNqkHTSJG2t
dX3bLS260oyVsxRJxYtEXAqfirVqgl3eFmUalQ5b+oMiFGYkdu9Dtqi2+nI/j7ozQKy+wVp57NHT
hFhxL9FliNrcsOEoJ5+uHMvHUjMkSTD5tOypgNg4Qr1GQWmOt1vWBuduIe0z6dOQ2F8ZOKkoCjtu
B8DgoFbc86WXIaVGfSpIoShH17qvhnIjaV/uJFD8npwtmISXZkl8IZa2Am7J8krSrLZvJSj44b0x
lBvsE7B7K98xnaMdfRkZagJXXvthS9B02NiLlobPtuYhaxwh/cv/duto8AVLDHJx46eO5CPBYucI
s15a4D6MzPshqpTfpjuv7TFyA49L9uImeBkyCLsfnWkE7BWvvHmmNzUfgp/xTgOsjX/mht2yu7+5
cK4Wx1pE7iYM88H2D2Dan0lN1UeMszaHHRX1RmEl5y8zYTMOIaMoZ08hyRIWdBo/BQLtuhFVdNbU
5rYKuag46hvGe3AaECrkT3lKizMaZfgxDXPW4AdcHcENsA6TxP4sF9TdgQ6I82HVHnzHkpAyl2IH
Vpb7uuKKFzkcuBU8xiHVmkbZAZ+W5N/cZJ+T66Xm+P7oQSBQ+Q0w7R9x04rri2gCHrRfmM4l9X5T
9UujzRfHIcvqG6TXz4FnT3RYsbTRyZifmrk4tk5VP780HgbDIgs0WG/7vG4aZt8pS0eG8Jmigx9f
SGAYTldiRSogPdfTb483MuOfp7EQ2cLeBwaARz/UYcDFWpoVqb3GmjNKZXcatZGxX7Yo3TTRF6yk
1t6hjNwwb/0v4gdBKdEqFLy11D48kWnU+bOQO8NHn0BHaEnmimFj/ED4pAdY4FMbOdaFjSh5XsED
vonPQSFtZ/SM470At3jMdWSbg5ClqhDY3KdxrAfn2OH2KqJKPxMRrqsalkH8ATxYwIsHPSyH4jYH
K+M81GsnExlN6DNOQhWPM+KNs4CL/rf04Me77h9/6fK8oXGf3N/svyK1iAcSSaFIFgBYhQwANVd8
ebtJOQXwXNeIE4rN35e6DtEEFAxYxq2J7LKSj2Qij6HVTAgBU7Rh69H85mwNmISgHb6pEatdHMer
urKG/uzso+6ND60gBEl/DrxTo6NJ9EZpW8lXpLg4/rkVSm4CunrIAIFfx/R4jKZE4TG/sb1Fe4wm
TqsOFjwRSzQYUfJ/ZPlF44jsSAIsUGwiBhFrXi/ToSG+3dXIS5E451Uz/5mor+3KIwou1ReVisCK
9XHazwTsr43yKW3WHaxtSNfEAzuJhyEFTtCEkn5FkkkcyBYP72Z2FYt+7dDno/ek8ZVnFBIdaEkd
2U1AYt0DhZf2+pPSVH+umXrkEboCPmFp2gFHRxHDLaS0Uu88zgP3ZxhdiDPRED7Yn0hp5Bv4Ov4f
3xSUrWg0i9+oXO1SoE+rfaCa4QI9MF7clj2G5SBMFSkZCJF1A8kjExu8I+Sj2henLeRNfwdYZyo8
GG0+WsQMM82vUUeBKW/wegNTH/sz9y8TrNLHpJOpKNFO6s7j9UV7CIMFLWZByG0tO9Pr9pyL/d6c
G/Jf5xJcblLamGoni6Zn9nvKMFthYEbkitxvhnTcyjtIBZ4ggKHvrXz/p1RM6lD8LEoWUp0WU/jF
RRWs+byZu7/pUNVVn+skbiMwb+JIP9PQLqT9GA6BJSkJLV+vESeGkzChvKWxmf8DpBB8y0Gh/CeA
5sTfyf83+oQzxb2pUpiSG3C8vTlh+2C8d7ZLOrVQjDCXP7UeaVXT/cIEqINXlT3r5n+qPx+Ad97f
5OGMZLwbooZ1vf+crg1Vntsb/fp//1RPwTLe6ttd3inFcdsOvkJxkQXVa75amuFFBkOzf55xIzaa
wCEiJM/wN14UdZ/ASEDk7tYWy+ORjcTT1avHw9XiebdPicqti1Ttpebi9RN53lDiRsccmLfvLwYh
2QvNH1mDtBUy5Uf2usygPjuxeF8NjQZmD02LLHFS9/6aB3XIJSe38euIHMYl1vVF/tw8Wgocai2L
4bWHmryVQDIFUnvvV9bSDUJHfbRVu6s1HfUHZaLd0XbQGV2iIjnNryuL9J+pGbaw8fiop5OrMnpc
WgYVwIneNaICBRMOWJtqgsW2HzK18JAN6ZvxNBZ6ZivuWz5uU88ZSwIzJfJ6yh9gVkGfDwdjdC+Z
OsAyE/NT/cdstYPiTeBYSVRKh5NbY8m67rdSIqzN7xkAmBmSvEeA5DqlnpoMhjKUlR8t8s9yjNgE
LBEKMShfpGqR1Wkvj0MUTEERqQDRDqCjj6eZVzYBxRHOI5/6diAM3MsgfjNzDFzsQ7LckKdcgih1
9SGJ2DjHE/1i7S10AlU82M3WRDjKZ48aNDqQ/T7IBAaGLcG81KTq7BthQprWfP5hQ6vOXE6aUf1m
5jG2u0B3mQt0zXJ+cut7pC5cyKxRFi1GKmK/nYF30xgo2Zbrh0fTVSYyndBqfKb+Ta1SOnqDttqI
hhwD5wkM+KLDsKisLE5NNLIPFUER9l1UB92hjo4152pEunkaWWTeqhCb/5ZH0JZWTo3zYqs/nJ0Z
taqRWo0TYDfs/MaCzEfgJUjesFzvioKinNeOQHAy//Gbf9YIT4xVuJXn3Ssxc15+mAepE5cm338f
CindROSDAPQD5JcvP/AZ9WhFcJJgl51bdi7ECrsfAXIL14k0VCQRZFpj0OXCatDT3luNgWgBsT+Q
bT1jFBvZrOX48abhXffdakrySjcu3ajpvgEhAoKuO7JJGpqswIWb6IwiQT1tT6gx6OOCqv4ynIR4
0vTHtCJHxtpa4+FjTpswKeOMqPAExBz/qfM1HHNds1AbTk/lrKmFmV+hJwtzypYXEs27OVH0Ib/x
7MvHL+JQvDmVNodwn0TBkFGoWIIxMwZdvJLQzKgt9bJdKDlLN+Nr1x9uroW+siJUalMBrKAh9OiR
/Ms2Q14ILRjesexCtr3e0o+fSWo00LakBqKwFhUuh9YLnxX2hsHsaClUKiVfl2F+rSyW0f+5qXJd
gm/+rvvYitdlXHkqAu8qscebaNzodbLGzXExjUNv9D4L5vbz8nbNfCswRvujh/OoLWCFvXUtnHQn
DrnDG6c3f2xlMvSOtgQt6DNYJKDCWgVbDmaAy3pz4FsSa7G5MCF8767DhMgjFlqkGsT8bzQjmUAG
fdL3DrOYE4T+o8mVdX0xRWDB5QV+Bj4exnP38htA1IEHdmnS5TeKHodWpwM6jBi/iAoBfJBTlCOP
MdMDmhVGUZfYjTtkN5ChW4/BPCZT6TwlXLW5E3mr6eWEVwYlnRTHsXbUx5RxW//lVSG8IFs2f/U1
JpiL73n7SjlujloZT9aZL7Ah6a/+mPz4r4x2Hql7QSbOqskECvGShrLjKXGYMENiZK57Z30ysYQS
beqgU2b5eXE1xj7wq3Tp0fbzn5VOQS2Azs8Zw4EPE/vmbla+uuMmb6BqFyKmK8AKEwMOnIiW/79b
JWwIzIhvVSH2qPlA8Q6uDqi5Rti81ZHycI3NZybz1/b1TBZOMRbW5+B0Ie87drp3n2BRL575FRxz
BsyUU3FnhqLQYo0o2ksKp87ftrEFFq7nIREf0F8FgPjPmMQjGGo9Bv2Fbw4Ha68HR7c++1zhKV0E
1m56Had54of+5rzBPJViSGbyhO+S7ZTuzvpzaeW7RSS3Y2towIH5pFwMZBAYvuMGe6QH8U2z3J1+
T0lBeK2ph3Ue7f6tR96QvNWmt4KQQiybSRU/5o2BgPKwzl9ISQXgAlxl/MjYbwMk00+hwd3bew2f
GS4KQmPL+G10C2V2iU9kBxej1Vi2ylESFzOQNrYhp9kIxUyptJtjCjwr6HmozFEApRuCJBQndSz9
LAuzRf+Df2Anv3zbpi+F8PrYr88rXbxtXPaSOkmpAhQGDaiPp7gbvIC7RVJk4DfD07TzL+GU+FGp
m5B68DvBYcFHaUg0Emrbu2dGs+IdQp+q3jfkovmAtyoyqodyGWrvhj4MfqAwvraL9vLuIAADOmB5
B1MaTqCX2zkv2E/3WcchP8Hds6qYjVLVgQ5mhX1XEA7mEZqyZnsXhx3X9KIcvKGDghyk2BaI86Be
F3HgtW2LfSfyHnWevoBTBiYGUSdUH25Km6eh2pHchUVBXfBQwukwvfitsoraoBRN/NT1rI44YE4x
Hy3IuwXUfoxghtbdUK1n7qycGa5Gl+I8jNrVIAd9cUs3EKLugAYBVavROzKOrwLwGKVn7uJwyVIm
dsB1vKcKt09wfhvpyzdm1Ibn/+EK6tDVIcFIE4u91Elj7LLlyrEeN9741/HxReMB1ZQnedZGgy1x
vNhy5iCwk1dKlO2zZ4YEacvaP393YIFkpiVZ/NvUzIJWnEsjBG1Qsnm/135rbw5+0FnLQRR1e4js
gLjWc6472L2n5x6hWZiarOv6RxVHR5GniQVy5xxZh9a2Ip9EdBA5j8f49UrkWbRBMSbpXFqkKVNw
Z/Cdfrchhsbq7MqcxO/Ce/l+g9gM8J0UCaOyH4BroyFUyPY5oQuDRl4jshWSN1BKH4KwpcHujOe9
3LgOAlZrX/Bjy5iovzFAGt6UTSDHZcVFE/BNHRKejO7m5IdBCFEXsVENK80QIzoWrfkIH7O3uRZe
aZeBYhvmwtYYpyGqzJs7nIKrU9XjX8ojS3b2XUZJZuCJ4JJATrlb8LwJcvipTeKiuYJzSRhHzzW0
iURuqPb5FAu2XLjvnJbRwr66JD/UOX+SX6ayRVp1aINrnxJ/ATBx3Ti3/V8ms2xAKzkNx75NDUFb
nbpp5H7HK8y7wuWDOnh+I6sbSnNrX/rrG6Sd9syGsx1JwE2OgwvzVzRJZxupVUyOyxbl4PDesmqs
SSV2oIiq4bq/zGG5cwXPO+Q21ij0xEvjP+Gp3ETFVfNyuakYoLZUMQWL9yur+m+WSTkQplWfUntg
SA+VVd6eJScydKK3OklQcgrpqQ7Sg+Eie+sK0Q2ES4xtIAx0LMHDC6w8H0h26aZwZ4eL8QBWrQhj
wA0uesv3MjQIwdC5efsdkiG2FUxuEeYXFVf7VBXipwutXc7ogQPuOXqboXeom9PXzWSLAM+LBtYx
w3tCylk7ZLKqF6WC0ci3JmRltKYCjEs9mDNkMbMA73cL+gmi+cslatOYPscDQHSjMisEzIeUVvw6
9BxZIkGL02ni/HMaCuu8/VxmLVJ60Q0JmngSxkFtGMzOt23Ds6G4Q8kQVTdFYCPQAcUnYNkxqVPN
wT8KX5EEUvasu5+BstpKxo7HITDLxLUrq6NMUQt3aut36udAlqbSkBi6ehXVxLi77mzvRjNmpP8U
eXzIux8+36hR6TmdBt9mYvEf5nRkjlISy6LM/gtHZfCVmBA36tzGucCdXxRyv6XS4XRlDm3E+3xb
+oyIcvdzCsmUrKgi6hamfsl+H1HLMtqsgWCt3eqVv/xjG04OHWfZk2DoWq9yuohg/OCi522C8Af6
9Iu9cIa7zG1RzSVephKgfCDUGo/MMlgBeXQ/9UJ7TzUv0NCNcYTpbbI5eabfyA7DiXN0LjKsKNLg
vxUQVmeOlXfNJ/bc48LZ8VQqfUPuftbScGpbfvb2faV7USRhogvQT1agwrqAEOuOseYAZt+vShiX
5sImG3205vGCU7aXjt8e+9gher4iM3Pi11yTRb0tl8MNs2rnFcyFscazW/cQoPLyOWZLd9Tzvv7o
lzHilA99UK1tJ3TB70yIaZ8bbRqB3h3Dorh4qNvin9+/tfFzpknjbo/8GyUy012j+l13es3MPeKi
+Qao0hY0IeZV/waKzMj6hMZ85/U1GFUNBwabakXMdIEPpQJYbFDQKFRxaFhQkS8qkGRm1iq92u0E
1jlJMGzRFqAbXsd3yEtNsqq0++4O4MSD4Lm6R2vnnXmJNvJfkxfKHYwGip4PeKDXQkcRxWO0+m+S
IzE9eGEsK3Gqqlrqdw76ByJKSXk/OoYKNWBVdK4v/IJ9D7XpmfHzHhTBG+cOKxrg5ywvbjj9hxot
e5FEoqSWynBt7r4SeBThK004gD01N7WRdiCvr42giNrtANmv22BcdZkL9cvBHaWYNDTsT70XgmxS
VikZhdMfPAcCkh5CBH4i+jqs9r7MYr81664drZEjgM4Wz5cHCStkeN/Sh5mGMTG1kNJrNJzKhDiT
0CxRz8+6tcJ1kLJ/pydLWMJkceXkp8+NA2wNrNdbGywxtqlf6kVMze1EBNLB2aC9nG4ASXFp0c77
OWy5PVKveAPwxq7P9k6V3hms0CohbXOKW25XotqcpREM3ZyMxl9OCLdl+wmgBmVy9/M20gcuqcgd
SztIpP5iT5teRvYPQetboCozPQsO3eis9YU7Hmhm2vYAJdP9f3Sl5OlBmN7jeXCkMLQdP3XfaJk7
Js/lAPsJ+AhYrYrKtUdT21ZyvbOkm4Tr3xGNwzNQy06ygmZK0vJtrjiDdqKjdGnGFxIiwxgCRk8I
jvvecIEnprI0JYheHtsTkT8NF9xV5DnrGesU0G8S5lzHA6y3qBdSZBYBl0afjRB6oVWEn3HXQWSo
E9+v087mbTkHoKLgWxNyTn/UFZFkbOv4KACleD4Iw5DDoqzksQZKDpHuyU8y/GWJq9s5wmW68jc+
sltWTlky/wriA90Guzd662Wr+VhXF30VekXW0a+4LIDUVc9YZu2yWjt12/y1/EAl4wggQavo50Wd
2vapLRx0pmZz6pCwO74v0NzArvKTBszJcEw2vnvSvyXftXD/S8pM1a96AHFrCQP5+1v1u4j65ACD
mN8efKk4jItBiaqtKu2dealcATEtb5PL+jwC8Mp75ddy5A8b7OGzNXBewAcyt+eYiSYVyVdHym0Y
XB+mvpbcTV+PtsgYZUylKIvqR6zZQKLeezDiBfnpRMfW7rlykgk85/DFGzWMYluwyS3G5mtNBSuf
cd8KZnwfbwRS2SUY5UYfThykglJaljFCEsx7ZhLyiMqC0rSjQGxUaC6QMSnWQyigeUYCy2fpeGVS
E4DOHoC7g7Cock02ATT7/U5IjL+7UzRRiFA5DtoIVZTaDgtEgVthyh1yTpEW3gFfm26KCotfM1P6
o0wM3vmHzZC6a8lWPrdPoWbnZM3IVKAMsTVrgGNY6l/8Gbb8PpCzOEfCkXPZqJ1agJ2S3zoXPY8b
GIbjVk81XfuqHi1+DeFJbhZ/iVfiuOPEMnGVz9z/4Z9c7DgCMYarWU4Cz3pEfSknElZYDuRTqj32
F5PW76GK9++ucZHfKqZtUi7C63xuyQa2N2QvBzlBtetgbAl/SVdII9dd7gQ+PRUkcphtq176cjbs
8C28T8qxeM6iWzVfUV5uTHC/DVzoL8niYpZdQ8Qu9FcQDrwnQ0w8sD2SCAvYTbQh01oW4NZq/JtR
FfLZNnJIV1nqueqeYF0OAkuF+XcoWc4OAj9FaJg3AjUAc87c/G8n7ZIZWGfmgkUeebgumqqNYaS8
gIwlHIOgYDdnGxlLTuLgpr04d5ksGVqzrdbtizNl6/blY14PIsnXLC6APTPPRahwa6soD63YXOKf
WEpbn/YY03NC4MpQY8X8vck+Kkdwz/sKrpBLxDBVfY/Wqgd7L8ogCYY692qmZsfgcdXIljJLlTns
jsWYGui6sI0YNo09eIZivfraHYQxMoPrT9eDWra0B1PXFZRYnIpEOhk2EDLvSnSKs6/CvzvOSB1H
OaEX6rh6H+bbnkkTLPIhUkBGNpM2uajeH/RW/b/LW/aUs9HFmdM1/Ziy0Bn8ewr6wi8i50RXwoEy
2mblYmnzuEcuEZY5DcMgeb4WOGGi3R8WuFLeS9SY3Jod59ZCbwkeLtSmHCHSIiUK5RmOlZ/Jsgw9
dvE7SzaJvTge+fFxLm6MlTdIN2AoOM5/u7yEVmWqy9+6S2bJGsoej4Lb6k+BUKXGh+8lkriX8Nyl
YVzRxi2tEMxJG+Io3ivqLFvXtD4Aw0s1NuqlLiurKKuvTwZpIOQyWKA/UGgnLYlAbjeVSyY2a3rz
SVRqfqYMCQ7f8slcsi+b2b+ey7zpf7T+BExQc+H1sobJJF9Pd+DYP5PoGbwMMeQIUqISk2H0DuEM
bmux5fNPwwTSSYicQACIWloyvpDTE5H41/Q7XuO20cxhuRtT9sUn+WfdDuI0NR6hhfWnLHpEWxS6
704CMAKQIFeBFOTr0jCKFpury313owrw3+7SHVQK88i8vAQ1w69mTpAJV2Taz575QN7Wu8j+BVq2
zpMFJ8NFwGgOrV3WBSq6dFdbtVqq8/SKG783pNotqQj7nbz9TMIelH+FJ2YnR6QiCDGiMlAL/wgX
SyZLhriywmI2SOWLrmWOapne30upGqqyqeisfDEFcjxJhiLzT5pF3gK0KIcXK8OlvDgYYQZ2wXYF
Zg1eXuj/9NDCU/9ueBlB9A5dgseUTwnNB3l0ZJdWIJnmvRheZ11UM/frt/ArwPm/4sFS4L5QBsCi
MwS6b5SybdI7qVupDESoM3EDREPGzTQwJJm9sQ4/n6XKunPcDJ1x8gB8Rds+dIbZbEPY/6DQAYWY
tCuyvlmbGd4mT14s5BQQZiBLA5BxVF8mehFY8alS2A7OelliPJpBwzk/CfTCGtOJe2B6gVSSQMO6
VOS0WUlw/0Ibr0NUetaFPSNPF7V4T2qd3PiC/vev/sIW3X/07RZSTntQKRvXqi/vIgfoctNL60+9
eOIbaj4H+zjItJ1rWT/0dwBkg3LmskQcSTu1eQ+uRAd6K78/kEWoGMBjzNGPcM7eSswnEBZHyyGT
a/Nk4FsJlOdd3XVhvq4Pe/J2xsq8qVhUpd1Nz4jMUzJCVoxfjMmeE0Lj2EzIIcjZs4mhC4SljkQF
KJpKJwHkX5WCWkf66nCCpITJbX8tJbFCoaWn7j/W5H87G9H6B6KVz62CQ66C7JxEpTTGjrbbS4C7
e5qEOUs8sZso3OBT+IsShH1NPSEYv+TL40KdCwV6T/YoyCcyMykyc4AtNduEHL5NjXL0rXTcnWgG
9m38iGXQyoVkL5VC6jaJN0sP0o/saaLaZSZddSNQkEfF6fWsxmNBe9ea2SY04/BV+PXlVoetrTPA
9Efk96Gil5ly8DjWnQs8EeHF5LhQn02QhBvMLZeZHuuyvC5Yta5M18Azt1DtHTsUe4oPimOeTUL3
az7Xyqt+LLkSkGJDK4BdgNeFEHXu0TG9tJB7iRMnx/pi6zkZG6dEOB4bHB65EfMBmoce1QrwmNKg
Bezm/7O6WWuKcJg77jpdYInMIWUVXcE3l8WoXfE1CoepYc1HQR1CbBQGXOtnwv9ujQ84xQZ5vw9+
ZD25vAsQdbKnyBlem2FYe0nNp1Biwh8cckDhEwfDB5YC/XMZ3xa1EXQTEmaN1SSSekSRn3qtsrL1
nRbke0L1a7LD55DOSK4mG2btiFugCLjdcFo7vGNFhYY1mmLrULcmRvFrF+TD3y2XAL+3A2k4wCGf
oXzs7HRzP25j6UTj0QjL6bA+AfKaXMIXwNa6aTDfdtb49OP4HzEFpNblN+A3L5XbSX15mu6uoXaL
9XvP12jmnOHO0hiIcDRO9VHbnX0s9nx/jxO10PFLSb3rg843nNrsSP1VdIj+b3CpPiiFYZqeeSUA
LGBO9Wtd53pBZrVjI8Xmwi0/Se2KqrYhMVfO4uSLkZ6ADjl/N7Qz0LV3rLu2c/BfMl+MzQO5QM6O
s8LlHObFr9/E+FBqCSpMLuIiP3ed3omZ+hvVcpwHTFFDXFGOJA9eUO5++Nm/3eB/vgJCRSG344vW
gNTWuWhI1igWsKEImMIyKLYgya47bYju7OGOFYc/D/5W5cTYLqdzk9u6pbJHlexE+tA4T8LBtSW7
kuHwrjHIs3ROukEKTHUVDkY7BWXkd7gMvYAOZJN5HOSBu6z98gFhA6Kivdi5OTF7OTLlS3NthbSp
NkTQ5MZELdqIZEHqm962XxA02J+eu5HY/8R/zXp8yl8JH2iq8F6swg+6v0TSBKrjhyZBbPnMgxsm
tkdye+2MkgWNu3db8GZtaa1JV+LUtju2kqoCN4dc0JLUzMveGUtHlb42UpBK15sj0ktNjsYwbVjJ
zE6IPZZe/3uMw/kPJJaffpaBwJGqj1QWTB06jL5zTa2qWyretsml5fEiDOPLAsCCAS8d796zz5UA
Y9BD8dEKKg5VEUbQOXLE1DIg9sArdWMSM8wVGTkEkSnBLgKXNlrW2Z0ni/qi/PeYQM4rWpUeSewc
O5PdJT+qoHo3+KJaqBDm4URb4c8VWATxVm+8I2T4OATLHCYPndKSmbJfoOgkfnXHSz9l6wBaWdYu
QqJreNsrk9x1p1LaJfdSicP5jLN5QlZZGD77t+9D4ev9djVW7zqzO/9m7khbxsj6qKe0RY6ij3PA
T2aMJrTM4lUmlxlSwxw25sMoVNFCW1Ikynn/aT8RS4oXlSv0uuZ4xzDzPgbMEQbA2pRwWLdJGJBA
k1s1oACkQ5x6+0aG4exln5WRodvpvSMTjSrRQil3d7p7wsrpae0tSPyNqdbawS2aj0i+4o+O8l/s
IndlV8RvUR+9/T3ufE35S3itUage3ACxn39x5g4lSk9WbZa8b1F/UCl83iJ33s0vpiFiicOu+HQ6
YIg5Y+EE/BZCbhlvWLxS20MysMEstsRvPNMz9ilO0yflwFAlhi1LSXiBODQ3SM863mubki0c7JYA
Tr/xrqs/UqfnDKGYbXyHZof9IqOrvsk2hUhsfgvACqKfWofc5kgJ6YPRA7YY2f/9SCuCAnLDt6R6
zwFFGEuqaypQnYzZe9ekmfrBvbmOMU86RbbXo+ueH5VnNUw/kCdqga8QMy2PKVR3xcMUbBWbRIel
HVZdqnLESO9IdB4fHMHUzy51q2EO6pgJx2DvLw/cJfYIEkjM4haHzwsaaNV+876aA1S9k8Y/Ztob
HwDuxHNs+vYi1PyVS2nxnHpMo6CMOmZMiSkYMGl59oysjbMmOQDfjWRuaHmv5qA6WomU9k0t7/Z/
MK9C0w5XmAS3EoI+CuSlbWu2sHcy9YEyIbKUHe65S7DX0SjKdLAMYN5nWdjzFkb1j56lO394GyrH
/zmhI2OyDO+fMsckueY/YLol23DaeKYAXpw/uTHuNQmC3tvJo7AMrqF+cVbHEwNoCaoH+OtEeV89
p3dYhYdI0w820PSRGmKHWdyXrAqKOZnlnTm/RBpqgisCPYj2Reo8Z5mdOodSN2lhjjhIG3r+6etS
StOO4BpINSh4FuCEgjml/l24fg2q/DdVFOjF41GRV75DyYoZHwduMuc2ZACm4l89eoqD/LPScG4a
fCfD2KIqETWClZKdj2EJPyvC1h4JrGobeEQN0n12003zLfZAKEBy0BpTOho/QmQWdlJ0HJ7zfGzD
AMpqjhaM2U+AsHTcNvgjTUVAdVZrhhyhWfmSiwB18DFkzkaiBRHrFQsBBU7KalAqyVy8rh2m5IFl
muUDqy+ESLV3H4bdEskN26gfWoATBq9C0PSsmrW1zcATO8SBXj3RvVtonoTHArSFyd/DEiFViy4s
UZncOO+clNfvLnoOCSOPkc8ifV6hyMaRVpYO/UAfp0qa8CqrRUdP6Hj8R9U9OcCIVq20f3+YlnqX
RAFeEfnEgNAoWFtjQV7h44HIZ0XG7COUhjiRJpuRZ2hkMXhpFp0y9vT/Bi0cJnVWtDywQaOn8g6Q
/gWrIuNfeqzsax/xGJKsmmt+YcgfeOiQrhe/48yy1a+JQOFF2m/V/Yq7EpBwxtdT5BalkK26Y8qR
mF/2f2oi3ipgXRN0VqEra5kOySmBgJHIpJYpJ6cT9jKimKONZFCPgJLBSpuNIjpjWO2QacOBkak7
lhovwnj+b8tv/03YGwiM+5d1hO2w7rWHrmWdCCDlywZx2MxNF11wkyMyuFu/5pR7S5YmjsZwpR5G
LjVq9ViWMkepjADPh+fKBqgXwL4ufwfsAnCp/XE3pYWyfRP7G/ZhQ2FpAHwSQ8X6FlECNG8sKieE
OjmJeRCLqTqJalrmih542F4XlzmnFUQCXoq0wf1TEiSufUW9p+2AFECX+e05ZnoFx82HJsevA5as
o0NCVi9L8VnF0xfljpbSWkr25VgKBKu4Bqy4sJdDA0TKidMXwnwBkkESro9I+ZrFYoYz9+rZbe2i
2T//gODAz/M9vnpSKBsOfMQqnQ+5dlAnBSJJ6kcbBuszLJt+247iHw/9c+f79p6iLN7g6H291ds5
c3suuw0Te6SAkj/w5N1z2/KSgb6QTqBtSr/xCdQKB1K45WYycwMl/82zt9VH4Hvk+oNJnRSGfjZL
EaVy7ZDgIJEW2uPQv0GzyF8qP2GfuRDo0K+IXgaibzrPQxZ6S3HOw6mo4Rf4kaharBy/I9woYLrj
WvsfOsPPnGm2F3a9qpPDN8OCjkQGaMgWptKqqOb004uoG+u+OJIrUQpCjZ1CRvGzokZ4qbL6XO8m
4epnbKRqbh36inwR1v+qytp/xjTdjT/NjAYl9+SCL5o6wAKycCQWiND8iHCml57icci15mUXWTQT
fLUItAi3tyAaM1KpWutx3LQ3RaLoRxKr817XezpdphEc2RiMHx5f+ide9Bq68ZxdONEJf9NKpnqy
iuvNGcQBuhW6mRaAw/ZtWGPzlR+LcD3e5ZtVVf0UELfmFvZIsEEyubXwjx91pggRvN0SPBi2d8jf
q8f9GRieR2szJYwMrctzPBK3s/kgH9dnU9l9ayMnHtanQBf6zfnmvMz3UJJp9f7bHCnD5i0yuS2q
khMzq9OBeZParqMoeog/YxFwiF+SdSzoDMLBHy9FaE9lZ9GDmLsnMhLO35j4DDD4aoq7zISV3AFQ
5MPN2K6ogJGuYULq4lpSRGQMuyUMd554UjeRvPqhWTY1EjFOZ8Mo+sN/v4NE7NEDbtl8C4mH2y4z
4GO+ab9gr0YAOONdvJ3BpKrFrxkDHH3GQWqJgcVlb4BunZvL5Ea6vOXYMm8Ry605iGgTDO3PpH7B
LxN1I4cgiPdiyeR1SGR0UuigqGM2HJLFGbQMrLdvl/S7txWT344aYaVBFUH+2SC2CWLJj3ZUxhtv
XpND+FRcawwRyJWcrfnaClVW1Yz3nQ/2lwBKA2DpyMWxob2boK+qnx1Z5TDSdaSKmlbJZ3v9K6eD
v0kM1NOEFJ5bqP6w6m3RoXZm0yFUfhR1p2EIMe08rqhYAGxVEk0lQMgXp8cPk39kuhkv/52a28Ef
gMVEL6CVRiVQxSOgez5MbWiRxKJk+5Z44xM7QR24Kq2m8YfPqEwcUzjIcjtpfsUTOsoDcv/qCx/Y
qU2JgYVhfrMgHPX+LeWY8LCKhbBbgHC9Cl9pGjBA4wbYrtvPDAVrZRzWsnouU4J6fiz4sKBEtGPH
GCpXs3HKeH4OLRQDZFhOcG+L4zDSS4fgK/ZeJksRO1tJKmfuN6NJU4BlMyOnIHb4UUyVmcm7P3pa
gh4amYi2QIiYkdkGyWQYGTy/2zBZImyu02r264Fn4T7EL/AjeQpqfLIAzNm2xi+VNQCkTr1cQDU1
0dBcxEOosFJLY9ultOA4TiQgzuzzhfrDE3BssvTHcBKATOrvuxY8fa6AQCGOcN+HuB5Fz/uW75sL
rOZY2ju7qT09pN09ibcFF6SO1wS/LhRcy/KzCxClUrXT03+8+yXt+6kmy3hBWzMCz00yhyZzz7MR
CXm0r1b6aXDb1DY3LnX60dAvpa+ZevQwPuIyAiGLv+smz9Zt0b40uuVaB9PhD6o9k9lhlVR+RJyV
u73TXn8LA2s4JV7Rr/pAi71ISyg26VnEjHXS3Y/lwFNujx0cSkWxdeXuEkTrp77Fe6ndBt+srfF8
EZu+P5pNnJfC72FTlk93NftIj6+fqXcKewpb6jfQwRhiIRma1QwpXv3p7XBlHaKD0vdGACzNXKZd
Jzpxe6PzarnpwnLgCokY3ayIwIqb3rL9cvtln/HqNzaDg7CgQjaO1Aadgnc9JIdW6/vuZWxjxYpD
A7Bmfa7rj7FSpq9qMPl4Z7NNUPnpnUNWr76rrNRGGUhzSdAx/Jeq4zwf9FHa7s9piN0RcExyPMxs
ZNvcHRwSzXB8yiiyZJJMAF59Lyeu8DqvY8iAgfeGD/NiZK8OMO9xYctuihlrYOHvZIsoFpQ3569i
Lhf9w48tgamfdFC02q5q4BsttJuZCLLW5rDf4RykPWuhV3Cwf2V/ZCjOEbsbUg3FzTjP8+973nT4
uBR3iw0QXMzsFa79uPsWa/EKqxxmc6zFhoIXaa6qcHmCsfrivVM93t02flmz6WI7FazA3mczBYea
aztxSyzD3qJzv1a9X95fajwk07lmBq2L3VsBhyuupAJL1Yi5o+YgBlaFRadhVm6O400MJbqSR3+q
HKPvml6+rxa0ymgSqlUKEL7rQUj/7Z5UepIGdpbE93VE7mvrsfroIlBSGGQtjbLFNjtunJPjQz78
pbg/yhq1NrqK8Eyz1qk5pClPhICytoerx7Ab+hpxWvGm84eTeZ0IhSkTMF3xfKLuTiO5doETSb3z
z/0QNUL8YpAMwxttlZsQxV0EuzfXIC3FDSOBFtnN2sAY+c0rlSx257tU1Igzm/Nreko2jhvCVlyP
a9bJ7STT4Gp3ETc2ZNp8tlLqZhSG80+yCajkbv4d6gvmKJ9Qy0leoEMMS4nyEGJoU2gMjD4b6+5L
jN/o/IzaDUiH4Z1QPRuc6dLxgnv9msvJ8FbTc+e6rojHjNxIw7mNad8lY9X5RqTSjlpzezRW19Ma
AOIe+hN2cerGiI5943ts7J2wpJGpDrXquHp/RKsxDigez3qjX2Zl+F5T2ggfXu9d+Kta7rqAybq7
CncLl4dEXzahGecEBWnUT1P/OzSBfU4fLk5NbSBTPurCPpB9C+GhNoo9PaG3JLFQsehOhZcFau/c
bA2g7FCMFAv7Hxk6do2a7XMSvmTJAsU63CG2HnFmkm9sRqiw3IUGJbjfM68DbqeRyRPhhjmlEI2M
oqBOp9G/ty/NHxuB34rSSwQYmfHbOFwIR+ayyqDtyjM9lJR9MBEUfRkWnozUc8u1/1219GLN5qdu
SDNBtzNia53o14ALWU9TIm2YGuEV3/8dVB0KLH3LKbNmCnLJKxSfv0wbEQc9d4uv2FgQH/gDn9Pi
HUMlud3tuk6Uf7gT/AGtckQbuDhkvh2HnBS9nXDsF9hbt4p6FswKH4tW8O587y7q2ovAX6p0ATu0
FQWLY2zdWGLGw0Qfg/zbrUdHocxNw6ZP6dZgGmYBfVr+UMIw51Iu46ZL2Sa5hIDo4N+mFs7YEFS2
R7XDnZ2WRpwepVGFVVRM9gJvGjE514qajTXwTK7RXpbpT8iiwg48VlOJc7/ysc2ma3CIXjLM9r+Q
gyZ/AuTfC0rKB4dGDmpovPWdwGkxMfSC8rNofh82kosF9OqrAKs9mFA5bgTdOGiUzL46BoJpYFGO
phsYdu4xzZcEnowEGPKeiaTs5gTt+E0C/ZyY0FteCmxsZLN8fZ82ytzCXEIvWjvxSAJSGNy+YIEq
Pl0ynSZrvHrN/NDOSjXognZqJ2CyLgnT8AMbEHPh2Sy2kosPCXVOTyxJdLhg44ytfOsfQ274FeZ7
mT2nSJ8sVrfItuJ4eCorLLA5Wnq8uYVoNSHQnAxCD53cBza8uLwIDDZBbs9GcgmgjTLboIm13kQ0
4YYJ/U14d+i7foD5wUl0EKlQnIKg/47m7rnHfnAiQC7hjgxfNfwjkZsvcGIh/IkdMZEYaScwUmsM
pK9X+d2z1LT9GtBd9KhMAZFnCFqZLIZExB7RMc2aGd1IjhYIWefC9JHhydlKlkXB2ZejREp4018P
JjXq/lLCwTop4MxifZtZUB7plc16DZ/Oa1HBVDrd13qSMkha21jyJmSHSnkeuk3z980aYlZgxpnA
XtjUhSJtg/0mOtiTfEs7nCBWN2oBD2XeqzPZYwKHy9ulYeKXa+hAK24MTIRDbH7Dj5XAesk64ku4
kkSrzwoFmXaRzCoed5bN6w35mMQAGHSfOGqqB0IhWQXov0N/ID7JGmcLWqU3Z+Dneqd21Zu8JIOZ
9diWWj5NFMjrpObb4+gXJJWelWT4+izyFRNh/JKAEE719IkI52GVgkM+GYiK15+CRJWZGbRdEWYK
UPTpFoUgXwmOWieeHgof7EZ4s/L7PuODcJ7+VpuwKIzMynorCDlUM0Fo18y3aLlExVTaw7dfiRsv
9DmZbJ6zAIxEu6BX7t20EqqnpbooqaXl8TBv3mC74dpHp3vjcACP6j6KGuEQSqJMselUmMDykbrs
56CHd/R36HLwNr3NSbOEg1ryRDNKN+KVGyuYfGlODWOWJuvLp3wiCqJNsVqstUsj4ZFfh3xWHQaX
f33Wk5slVMEsRqqjbX/e0m+48C7TAowu3/xE2q4HsX1hBfT5DfgMQazuPV90xU6Kdok51asEG015
syFC2A2t40F3EfCSNq1KuYPUpMZ9/FnkyqOeWZV3vPh7fW3REcFDpaVE+75I5V/muYqnqA7QWCL/
6wqJvtY6D86TAv8jdPLqj/pZe0Zz/5ROuVN988iCVE0Y/cbezi7Q7Fdnx9DgYYlvq4JLxXwYAj5z
e5Wc0qxy4g6Mvel24ax3Y5DiREBGzsbfsBEUdp7f3HhJh83r1hDkGkp7/KjLdJTFBXYrtA2EhyCe
DTG8fnhbEsNvzVTBp1qhMGKGwvLwwGdiXSnKGTVrEAJv+t9zXe+LIK9LPF9OUwl2Q7YbEEPsR0N2
FW5M8xjSd1ZHfKfOUQ0W2gAOHVkhCyTSaGxGVM+wwuLM5sE3H9ViZSKgW3m29FeSl8EaW8SHQcdv
706WNBaKlqOIIgZ3Yd4wkB3KuJQH/avXXwffAPYV18rs6eyBXFMz55pqIcE8HaXxABMNdkODDDZK
QYEWa/jlp5/5gXJLkHw1jZWYa/MFLkan6ScDarOzBDYwrxKiAeJRZ3BXxSqypryajZAiCZ61rqdd
wqPNt3bCdt6fk0p/lIQFA3ZzkYrAfCUKGdMYMQQMGBLILeiOYG5nvuaji1/ARV3+WRoT+5G7HyPS
t+OPoeCXEYOK6HUfkF6vaYkT/StpHODLNS/Z1FXwTpzzar6RR5C/LvZWurTE78+1+FXzxW8LsGq/
Je7t1HXX3NSv3MNvbgUel+YclRNw5bodQiJiq8Bmn0S8wtJ7wThCdnN4rzAwuLWup9D8VAG8uQxf
6U+v5BcPeSVjwvx5K+Llkne562uU7I3jq/7Mjmfq1uOCSxbZ2nOjGZyIG5LctdHjvtWzpxDhqSw6
sODN6EtMBssQiWXH9GVEp5LtXA4Gsoi3dYhQkJplxxBnsjOYz9US52YIP1aES5vTPx1HU/qIUss8
LwR8UgJn1XGEYEuFVWgO2ItMZANH9eZaLHwT+DHccHXBNXCASRdBjT9Y6JMxIeEpt/LYa0yqKuw+
fMbnX5p1ttr8/j1KCuZi2COpf97gH89bL3XtTAaVr7dOY+0owBtpVzATc/SOe16zZcAsYTd0Q2Ti
ra4d5fl3lsEuA1ZKRdOBjCSUDCN4yd2WkG6r69Ce5dG/dBJ7+fpKc1tIOymWnofCM/L116si/cj/
rWU3DjIP/BGG6ITY5iPSzo98Dda4jVYAAOWtdRowzyRS4qrJHsRV1SExu8tR8QKhzykRksYmISeX
lHQTOybOrBKXOlhi8o0DvcqCZmEnGv7a101Q3Iw2ZR0JEQPvpGCBpGwlq3ISlEbqOtODNaWzGcvf
4XLJAk2B5Jhvg3Ui3lEG1J1RHJhjR2JQvMhwz4hTLgX4qEs9bolB5v/BvKkwrL8ygbh2lHmSDiUf
NeHUqLbQAIRWMRUtk1pMpr0R1UXZTOXh/qt5A60QnutBIftBQ/8DT1Y4cIz1jDEUixShjsDSkW99
rmFqryjgxWWlzpEARjzvqymfA80mSe+i0yOxhq//05O+QXa4a4tpzw3A9m2M35PK2Jt0jZ07ftv/
3XIm7nKjCFiklCXnGb7YVJ04HormeX9Q2PNQIyjzWvwmF9kPb/aOLxrgqHjUYT7FLT6MJyLc9jWa
IOTm9RyndeDZIPVNSOhf1UVkCtCItdqa4Mmn8c/IxYX7P7FRdQR/NVri10f/OUZ78rrj8KCqHRUW
mbRScnl7eyEvOKGfM6WKxaBMn6YECzlVcKoYjp6ySr9Pcv6dVvHu+pzmHEJuSWKXhv0MmOxlliV8
yAza52lD+MREy125D4bem2+/gA8+wtMgRz27N6c64Tbryksqj8xTxSe6Ah+ZcUVaJ3dU4Wy5xHM8
HEf2GCWUV51UfKrKc+bR+E5VwTuqBgdx6ldRjR1B4wbD/U7Wwe3o2L0S49teg5sWKv426lZ/qWOn
bj0BpKjUv3LaeiJnLFs3csjxOgwGYSjQ0aGq3sZ8mDnaDQPuY+3W083xCNCDlLIxyz2GmIx6cSrD
lti7uwut0TclTtCkBwwFQpus/gCpQ0YY08Fo5F8PXIlkoJDB2NLgMxmW2zCsVCpeOXuqZSeQ+Emx
ETp+vuynKo7wTQLNhhJ0BJY/JQJXZTAG/U/hLqp3hRQLTFO246NB9WO9b4V/woglt9GQxI07o8CI
DnAH9d2FOpzRTbSeSOpZa/z/C48rMmTwOoLya1skFGSOEC/lK+rr8YDBOCo/6K82J7ZwIAd/ppif
c2NcxRVGLYO/IwQ5hfv5Gtr1Y1FBXO7kDsf2dhLJ59tu1H5tVqYFs8AV6ri34PcZ4NmKIO7izCdN
MtyvG865LEaeRyrcskm/jAKmrPdWMB0XqREkEqJMvBeVaNPaxkJ+xdv+JEMPAYZHE57Vf2s8xWwj
up0Swp/3CIYfeyeba++zTNsOgBPXgZexYiVPFPMG8gHT9GyPDk4CmqW21EyIF6EObMQvF7rib7Ri
V5CrurN8VGXRTdPha1ieA6Y0IXw+cmL9OZBjmfMQ9jfeVOngM3Sbl4T2jmsbMdTle+b/EWkVh6+c
X8+b31mlk5HrnVVGYq+ZusCiwYFrd1SQXo+L0B3SzlXGtY07hGNYbY8VJrGVSf54NORHMoGzQ989
MKMcBXBiGDerOKolL2G4msNDwfA+HLuacF4H3B9gFH1Q2zTWiI4CQ+cyzf7F95QkHl0dkcN72Mc2
IBpuFili8znr3r6WgWPT555T2IBt5kGIVhenb2o6xZM9qM0LaWwlafONtTH4YhQnSXyeHuQhL9GM
VVkbbeQzVcDLTB0J9LpXOntKQ2cja2P3uSyNmb2l00emqNJpeU440YY14UfXfAckOqDRWTdggHyY
2LkFiIylyKqlnKIyGtpojqqwYVOpogaXEFkT+KUO0K4Vf7B4wA12dz5OSebDkpq28p1E9oLdhc3n
0xlFIq7p/rannx4SJh8ABMlEs4Yi+7keaXwYVFvAEr6hgWKPbEwe+aKRoMbnCYsj9gYH5sZ/DNAf
r34cFt/cAInLjVNvcIcXae90kUhtfefILoBXGVpEiwQd+N2WU4J6x4XMZAo79kcIfthsIhlYjD/a
SJqsNetV3OH+9eKHOxQT0W0EtEimdQusuMiJtkCJf2S3pzjEFCzWN0kA09ShAEqQVKufkLwm+Ttv
VJbsKRrv8GQI3QAj78V8piQvKjI62lkQTepRcnyUvnN6oMLatARAuTEL+RNkUhDnnh9PlB2WZS40
etzHi7+qgpzEYa8SYoggsQL1FZH1bmeAO80tkNMX8tKKp03ac8itUg9LlL+hbFCodkrwpyGKBtzM
YLmOLU90hcWQ0XJPnXI1XBBGbdQcLl7ItQpRvrWws+q6cNOgjhTT7G6Lg2QnhEpcIm1G6QGZ2xvx
DrXsjS2l36p0U8oTtz+ou+kElXTcizC1z8UZZVAkfcAj98LaZ5O25iV3VHjG6vNyaTX9Pv63KEve
3x5EUFz/5JCp7Qk5/wy6U7xd3ofXFJvQUmCHFUklnIsnQPg6WnUGmRvADoTOUaeFSY9W32bV14uc
qkIc3LnCS3tVhcVx/a8+Mxn29voqxVxiUMeKuYLKhzyy7/IkZWMyxvcrR5krQKjflYxFOFPz0iUK
b0iBC9coHvAjZLdm6+H/RcV7zB6dZscfNw2H1nm+GqKOkncZ3dS4ezQyoM4SAkLSe8ir93VH63MH
kkJ4Bjttq2ec1MAgsdItphaqdy0TUWNE+zKgPGXWIcfwqcX3Oa4+r7nbgV7h4ioz7FyLzKdF+Vc0
c7gDRD707fJ770DJCteI1jynPWcKFpHKz3i63GndMjdvaBdkax5lFpFvZhyjGPI9RD+U1VihwFE7
9/NJrvOs4OFB/ZeWtPANWn25eJq4gQ6Jeya3ywzFbtZ7bEr3Oflj3DJEpQQYj1/1nwdBT9k6VcvN
4m72N8rklJ633DnQkIfLdH42UG0CXqYxw2S7zQZ+cUyPCfOjDbsGCSNxPOsv9wAyHri1A6okfK+R
JsBwOW50L4vw8+V1omBWweaBo3xJjPkdcf3juzezvWls4B/HO8K+3jNwdCoOiL0OPiE8LT5WxZiQ
Wcw3Z7AZ6lQA3PYrvIVZRc8nynUGSbey1q8RmNZ4QvOW4FP59ifH2+sHYTpgx/8tphNuG/w2Ju2g
BSSG4HTT1BqKfgRTy4KLdHE7pJ2XeQmNs4IDEih9MlfCrxbUKfA1bkg6IOs2m5LzV52BdSp0s85x
SmDpx2D1Az5NmdgSMUEcMGJchhIhRmcLX+UXPm0bZ+GM+f4wdguDLxodTd90Nsu8v7tuTX0ZWeeo
iWHDYwG/pDMy2U5uoKmbWlQci4of52NFTV8nInBwDVHEI2OsEYoxqNb5sPbZoecs9sOUzwXwuxpY
5HBQgQnNGZt1blxhlXo8L9rA+EBH1Rf0ZZKAnBvubBBsXgxp022d66xtq0I0CVL0KzXOZNdbEfYw
uzdnsSu0MBW2bz1JO6RiNk7UG7G3n00ZxbIcKTQpPmSbL3kjJTX1lZ2eosBw1AfbpfiON0RYRD6D
VNubBYGGVq8wl2247of0ItrGlKGn+SHLSTZiWOVUuLdWOmGICkW1LZDWnLE+GaTXLgo6e4eFeMXl
K6jgYwBh1gmMjXQKpUf6I0eZbrRTG9VgSO+GAgH9Ntbvsw7CeaQ4Qzo+fT3qDIit0uZw6SlqqA/e
MDHFcNJZWYiGsBmY3Kylwt3Ei0qwT3fSRtMLVuMgon0BHM3YRL3R9RAyLzO//QiQ+d+ioXnmH91A
w6hEzUZCK1yEGeMJ+sR3O0wHgRHoZ55Iy90RUNKeMpU4j0CgxmFDBVpAej/7TSnDWzauz1/DIZJA
pvPBBwdPCffSJVAnZNnhmccHlEp0JRWTKwa6+Q3j+hKvbhpFMvXFI24LjU4R8yCxOL/h5Kakf397
hUq3KYTfWRtsiOoA4VKTHpMCl5IKhIIt/ZsoKJ/3eSOULpsLe266F1BzBicBDScJk6a8fSKxs+Mj
7wsrpd+z7Kkm9DOr3b1biVPS84uJryIZzhVtS2MyZqu0/Fu7VOgT52HVIwdqxGEhXN6BOotCdlPP
rpnqVdYwEXcKrKOOIntdhdvEydxbBnR7MW9SPzK2j5ZG3wq2Uz+9A/FBqiHaesRZjp1hINaN6+gb
S3IBbl2eds0j6aGgK5FWTz/hXk/qWNCMVacety8lkiYnNSjUrn3Y56dzYGFjH6vxYTnpvB9KDyAB
EkqFzbkcFB+14x1n234ZAHaEBheGVuTjfA/pi1uM3mVzKCfU+BblZYtsp28XwJ9v8RXmlD0cdTFV
+5X6SnPkIjsdOvLwlffgDApnoEIoVqoh4OPQ6IYz32KQEcNdAmJySzPfjILFOhIZgKhiL3wEteWX
rdMnTTA90+i9Mfu854CHzORmgrruFTyOd0jH2swVb8uKr7Zt/8zwavjNVUkdR4faXszrGTPRhtia
r6X5PzMHse7PSfbR7wQ4TT99ZTYFQkcumTaaeWLm1wknTZLRih9QjxGWvM+JTtVf/FiHNou68Uge
++UKcl3cjrRyAOt6IU8pJIg8wnTHaki51FBByTTPqtOh7VK+yAGkAgLIh18nFC/yKzG1rYHkZuvA
l5VGJsJMQ8wMjkBT26nQPzO6P5oyu30zkwzgOB8POClpzdlIGfNLkXllTvRumPgGzGGb9Q2FRB0c
zdnTNz0oCFFjLh8O4PKQGrN+b+UhACfA7y+W+uGIq3Ivdov5/F4VUYWUHylwDPqB1/6o5PdJb+vJ
jWrGxO5fDyDUgpS2totkhnmL36wP5e04QNzrk3vyydj3VpqD+OBDec3EyClS8eggY1qKRkb+Liqv
jgVOFISKxwAccs+sSvmw8T5z1Vx4ugw2+244f8YsrfsSkxh201+xTsKGMWUo4z2AHL9ggwxc9aFL
cSiFMt1jhOfoRuxtzxII8QO8wfluYaVi0hvQXP02No4CGM3qhnYxcmLdqoQZRDjfnMOqWzmGFGBs
wA8d5Wf+R1clOfzusNbfgXk+nNvvKk3FL+Q0+Ge1fD8wk0P3GNk366iNHpd2oj3xvtDYSEIBmO8Q
ql4tBoHbJOvM0Qix70x8A+Tc/3LgIJU0jvHh0YHqmYprD54UDd7XwwFElwpGhZr6CV5cClmdS4Yw
VO+nmA8Ien7e73tUdnB34e5cXAH54dipGM02+jzGvYfV/dSrDfYK/DicnheoYOivXIcFh15Ru3Y5
c7yGk/Xn9cPgtlPNknRCq4JcgH52NkEGz4b1D1/6q8rQk6OimM3dcCkG/oDj46e9c1YxzCRCnP/C
oZpmWiyDHGBwvg/IL8NCj3bQArvewtZqxYzBH7FACVIFJptUHZVupxSiWOgdWdNma74joaUym+4N
aGaV0WmUNnxoG9Z2oBAa8zlb5iKCct2EDc7uoyZnzrX8T1ocELEsvgIbj0iUdZcTsJRHH3dGYlZV
sYW3UY3DDu67PJUMnCV/kcU9tMa1o9HPuG79/6jcbgjDmK7i4fx2Iz01T9YyqxAsukod1aUvdJQV
rlb0ES1yUBf0dvdvagIAUgxSuv4mHaOyXzkK9xCaWoiV9BlrYKn+eZvRWNaMZi96EAs0JyTT/LoX
HAMDWKOE1ZMJSClZVWtMeP/ayH4SUlgYJpdVfWEFBthbAOzf/8YCC5b8lDaoc+CvQUbclmwUG+6Z
PkeqjhzWUZzyYlMbIIPQf8fHUfTwBfypIFFLtUWvy9ES8QY0v8k1EdQTOSpN6hi+D25FUqyTLGaw
2v4rVcNewJcs+Hdj0JpKCBIK+xCHIL8FwWdkvePTiBJCC39ptz/9PBjIYeMpmtOHGuQmGxRLNGPX
bw0oCgtvXSPVM2gOYA9FEjrf2tSALnCxa1f1GPF+m50zw19TUMP9zaqNqY65zkPkoax1gL9t2VNL
RXm/etXv4IrJD6ZcFxn7UiDuiDTrtgYs4sjSqyJfW9EGo/TsXVA6ksIKIzrkWbRbVrG1phJnGbVL
NdQNQGGjFhFk3ae/ZabLGMJ3xqB3OzwuXWkhORx8V/whCWZRiHMZtJ9JouufN1aZ6SK22FwCsQgz
bVO9tI9mI4raIQFP1m9bRJAr39RMGMM3JkgQkE575N7v2rTsZsW3BQA2885+k0vLo1l+vhP/CnTs
OKWK8AqIBBThVGGVg/rgYYxtlKVox2P5nN1NG2gm1B59wIjHsJDw6vZciUzGuFf0jNvrQca6KPk7
44CYtBYaugoXKcQVqtwlg3DiwpGAheO6TGbZ9GAswL8TVGgQLKzEZrVtdpgQMyT/HL/2hYJxZF/q
+bbhIXWUHbY/OZbcvE6ap3H6oGBYjGH6R4swgDF6EA0U8owh/txUGHObJsuzVje//IWRUdBj69SU
60Giu7wfG50+qvTMbufD8+KNUnIJ9lfuA16UbJNaWUdL3RmBCThi5Vp8KWTw89gQ+Bib/Ci0EzHe
0i4tIrq12HL8Zui8l7x3EB158METIk/4UehWJtj+k19D4ZFqGPkORoQpomXIoLNdxNotUMW75hry
ZnOa4mS09up2vOS4BxBYnjVfAtwz0qo6of0OxNApjhG5BA9jy6LRd4C/f5ZVtZ6lwsJ7HW/Dgtzl
/Yl02psnM4OrI0I1gPVJS8igFORMRMFKAUUlFr9eIc30rRtblYeZRf5nV7RbmDCCf5KLwEOnsNOI
pfJP1cd4iQqHjw3PUcYRqtySAb4ogvOlS2NsVCjFDbsgmdNE25z/6m1rv0vfUlqvSMpWRdoLPRia
Z9wsjPVY7fYBbLT8wVvGiXeJF1G41YRdWnho8uUCUpYYNy7GV1jh7x1ay+JaYtfZ0IEYbz4xHODT
q4u67RO9jnsTO/uqixT1ij2UjKdlHhToWqQGv8OPDWBShvfZyeBoboHpY4Q5w2QYNZGJbXt7yhhR
JnXM5QkDqi2vERgg5mgLw+O2AltJNAn5o0VI/Opzo+h+I+L9SJJzk1VNCabqW/rYjz4ToibEWzBh
fNEQ6F0ljfBRdVKPnIQamoJ4eD/OQfUbJhY2o45faMwr+Wv1DWlM02AZLZL/eYbpu2gNIvSbUcFz
jJY2QDoFabXDQtAqxvxzxfBmJCn6EQ72hxEEKGroN6BqthMYGRigrsm+TWjviqD/+/Jk9kU7TY5U
OdnGSfMcAl+D1mUbvHNE3AaN2l+iwuiJEw+WSqCIcHb1C6U0Y9jZlz8Df0RYcEFPvOGp3JaRuib/
T6ZrhyJCgc1mqEsvn2VoamxPdN9a17vyDQwN+bpK+CzIPXGlgclWxkS6ondFnfKmiTJoFv1W67Oj
RfyeEbGcfgUCtTSgjo+4V22c/OePotzrF+FGOwsmN7lY/oLxqunPzl+ltRH02XyEpCHsqI8L1qau
NdZz6WbPVwp4FpxvYzqazM4AhcGRK9DV6itj3HXyLWMvO1Fn8haRZ3bISQFArw7bejsKgQ7XKg3k
mPPwVW7KsMrd/zRBvK+dwxSZc8+WkL5VYzUlND5ShoLKEBapYaTsYtfSvjYIUL3Kp5Vp0FlmBQQ4
Mz6fARzIqTe4nCBNDckwZEbnAly49xHmGZhSWRss7kkselAtkr2eLrfkojK/CMdhlwZPv7MpImOx
to7WzC9q1iS93c1gjd6BA4gK3qYPUt3ee1TY73FmFZiKgPa6lupNrx4e3xODPc9NyLDWaDrBRZk9
LIpRWgOZOLOFnNtNohL6B1aD6Pmpc1MzT3nX7haP/63iodFynL984whOcjoAxTDkUKgnUG9fcZjP
GzflXhPat2Tgw2b1GFs0Z05wFGS0/zMgVyYgydNslQMWW5MtmrS1qaw948ktiusgd+5MsaQAS5jO
XVxCThcav6D0IN6SA6Axg+X7pidAhfzSUdFq2DVrmfWrEBBvFQMN5vEIcOGWbaE5cfPIrc6gweY/
/rVoELQ6nePMBKlzD3P0R4ogPJno4OTiGSIMN6bh335/L6A57hJ5vNPURKVrGMUxDwnA5egkhAHL
JtKdBu29sKpDEOVKaV/ppc63/2wM7HpY+WNbmBAfqKLqBAIub6iinRflZlvsvOk+F1UIH0eVk/ES
Jav8oBM/jHwV0r0qDRxj/dL2XZne5lbdAbsqNpXTh22rLlhck/3ANUVtsoHzqQKYIoPoZWPt7mks
UyHUeGVtGGrhi6tziyaWBViRUMXt+I3u6plLgusRo7BDARaN4nkhaxfrxxquUufF2UUtqgKmoo3K
pUkVPDaMl0A2MHY8LzQo3HHzcSQy2XoAvkABQSdy1I6qKuYtzEnl34T2M/SkphFpw/Hc5oKdGwjA
qTP4lR1WJn8GPAFihoEQfqG+75Lbjjk4v3i9Te+bi3yfs91V9c6mxK7Ako/M0QxfhsKFoGM7607D
gBmQ5owIrB6vRix3VuPHRrVhfQIFrOKg05O9RnFLflsgDBhbzNRdrGu8sQbC0wCcMdUFcGxc2k0i
DCDW2cMXo2B5lcsZkqeYpuNq6cv58kCmSVfpth32YnDBHwNM+V++Hqy6AqhA0urH0FZcceC3ZIc6
GIh09ILwB1JP++G7kwRC7t09Cotd2EPna+wcXhiWGj1rvaHJJKbwI3IaqVuwe9rW4vAHMoh6JdAo
1ClhQCxUJO6pTty3wudttpadPYG6TA3s1edVMVOI76aum5jsVG+ZrdmLuGDHhqjR5B4QCHXVD54D
0gZgImoBU40/I5aJDP8jcFgg7NkA71nveUno3pa6F8DmC9caNKf8DvMxw+J957ZF9Wtp5Aq5iTNr
txqfiOE9eUg6eR35V16f+rSiRn97pltZG+PHlm/fD1m/Tn9odvUoG1w7UOw1K+ws61wxDF4c1qnt
DnTnQY/d5efRmKMaeOSD+eEESg41yUOTrtkjxcesLhcTxUX4SlE7PE64GHzFuFMVXurIWvHUqfOH
0V7PwxXyCPc1Io4kFHv5zmy1GpO4Vd40U5FFOG/nnzSWprwBolpKI+KqeSmWFfXMyI8ZDpuMry2D
ju+45i9EFmuGaTGFtnPjUBCae0dgb+UhGKtbhVumoBMkCmVFU6G4XR2G8q8HOhuPDVqq2qh04Rfn
GtV6rhgTwW6aKVNU7PcUaAtKNzvl63igtjI23XAnYUuCh+Fy8KGYcWWYpbx10ZVo0jxLk1+ji1mV
VkjQHPzK9nCA4V7aeb7QdW315weJ6fB+51wx/svw5CZe8vY64qNkNju98nOUHNMrK/5Fqbii8+hD
/MUVUuAOFCIgUMedQPT/yMr8z+AzhS83wQEKrWpWmtJZiZJVsWMJ9TcalQq+NFWl7eeZUfKNaUHw
ggSYtXeu+jaXT+oBVJx3eDjk3q0Ebr6uznxTL7qD76uw2QUZXGn0nSQkevb9Pe6xn3yZI46RRlX3
TTWnyw/437JckejM0NkNEKowdpmYlNjksgnEbeI27tBbpkNZ/9ikLWvTjXvj387sISOotJ1N8i86
hGUQed1EuWTFxD/Kh2y9WFxcq+5Qpm4kEMOX8w5f9iVgGgV/GB2zyO87ij7yfC40rC7GE1bY5V5g
J9dCBOUPr16rJx46jWgR331V6kTQnVwRAVSyLCswpdb0MmMkgWOeBGN0Iq0Xl6kTJ793QCCBmGuU
+E8XSP85UnzVOyeapJmsiptru7cPdlZ15FZmHVsKt3yEakodTClGEeNjUroAzNG7yZukd4gZk/+9
PfzPpAC59zO/gYANZ52kyH26mKth38NL+aSn1aSO+MjEfoRn1w1JFvIeX97MNNx3Zs0YIvNNoP4V
Eli7PS0kXmc9wXPVn03+/cVpX76kQDKd/lSqV33P1S4GXOa9dWN5m9AHuy/kmKSOiyl4hIopzG+y
3B0ciSYE+uIQzDfLJOCBefZUmwmv/xImSE/2mplSTjVF7NdIm+MaDD90FcvmhRmomT0NX3IbYhEr
Qeae7QSwOscQOPq9WvVqfN6/DVrg/A6rD7b3m4pf8HMypsCI1T5lObWNtTVHQqqU/wjEDBDM55sD
2sjPfW2DKcs+O2gUjIIYpD+vp9pHd+joeD5NDba7VWJbOQUIE2+5mLUUpJnizH3ja3oUqqoMvuwU
Y61G3NaV6ea1QNNTS8Kd5Z2t2OJvq9UX9tL7PUUdRH4G/sjOYcljP1XtL6t7waOXebL6jKfiI30p
tfa7DgbVwXQw0hPUvuT23s0Kk2rSwUMVclMSBDG2GwabWKKMFsGf1kuCsFMI5nNAf+QEL9SoaL73
d7GJrQpfq2x+hozjJdOPUQ0sJPTqxw4pyP2CgmfTVQ3r6A/sAzvnrfWvM4t1zNRdxcoSdkkIq4m6
YeJ0vkY0eOP3YnI2Gh63ewIqfmcp1yiuRV9+jJrGV95lmSWEkcfmKN+y4bkTHn0VrnkTe9fdTAht
5btOWfiIoe3/WN3Hm25rw54adiEYfODHtFmMyCTXCrjnbH/PjkU0Z6+ZaV9pTd71w1rovAyrntjd
X/qbixOB0H1rqNaO3i/6wg7bCUun9tUfAWVowQOmjvcZ7nnTxoqovIqD2Tuj6GkrpV7+1q9HgQBJ
y1lVdEjY5VQkfkkOcVB/SPBC4rtOhm61W9E7FyB9Wccr0k2KRx/847MubW3B/lpxjWQVviMkWN76
p8VWjqHP6Tha14ByNNU1j69Qb6oA4Nqp+nOc6nHj52zlqYUZnsnxmcoCOI9gbKOcgs0wrr4O3aLQ
V/GEN0fUNVclFEfTGd2zX1Q5TVoq6q5Gk53PpK2xZ/4K4KyuCYiXjixC7lYcpFBUKNS1G6rCpTtA
viq3RiOj/KtxP3KyOwEyTr0blfq5F2nBKYOZwaMpig+gacFYD1+1D+XEXPFbW4PyMYQVt9GvPRou
ME8IYUELUIvqEgQU0GSnF/JAbLt28NA1u/lO4ZIfc+GS7zmzw6OPDIAkn0HcFVnif/aOszMJQqzy
RSbnUCQyoCjVqxejbSNnn0tHa1ew2CaLCQnyv6QTqcxoxXtGjsA7MXw8iSKUNyP9EawtbNekGrtl
rnQiO8A419tbUxKmbZZAt43WyMlU5AyqJg7f+n/Y8gUzBx9JArEgi/XJFfPfnlhdVR3wk7EEiXZc
sBBt3Q5X9G01rcffJWlqQJhxKYYu+BSr85sbiMpMGB+6zBl0omMeMEzmmxkqTjIlsQlXo3rY2eEb
tWDM96sG7NBqoxDbAfFZ3mlqsav3ANU5jaNBJjn/qWmwgvTxUkTcviKQrp+XdXXfvDFNpQyFccTl
MXUkFXL+Esar6/k2PeKHmY580pnCtFCm/GgT+XgUDBC9EvDQYd3dg4E2wfvevFtYJ5hvKtaMgGVb
Koz1Wt5wRE/k62kk2cqhXgJDS6utfRKgf9vZMqE4eq8N1Ig4czae787nLj5rC2NvbFtzos+ZKT42
SJ+WcnsUOgIxDrvgI3IlYl8zQj6Yv7uLvnzg/5iROkgv4y1scuTM0qZLvVu/9g7UHa25UoCzA6L1
NP76Zw31ZZnTjNLLOfGVldFOfKErRskVyzz+kkx8aE81L0Tyw/X709Ugcmni+hXt1rM1nmLMJxgm
THg5/Z/A3Uh1p1Tzg7J2WVQ5Zib8D8f01KtpU9F+XChpPplOtWaRYllQz/W9wGob7hN/YBOHPFXd
hvg3osCTom+g6WsBDhtfLTOibaGxL2wvtDTXd+hB4IUUNH1Ihju6X4w574z2xUWousWXqKRup2fW
IqJ/jAUX8ZdUbnKnACrQ78rzSEFzRG6YmqbS/pm0sLIbxXO+BD8WBRO85nKJ3FE6Eijbq+160jmW
QHv2Nan9aDUNP3/pvekHLXz6nlbUeNhWseg5S+UPyCmYMz5ozuIv0eBlIl3t03NWw2eKPruStx4f
OSujOMrjMvYwgGyixJf9QgvhFT68060RgNSqE16mY93AlL4OFxOACZFAGNsXp1seFLLWUR910fFf
Dew1ag4auOjVss2QyRjwv0CJD9boc9OrTTVmt4KkkSkU1moL8T4w5mAHyV9Nbambft7U4mzvEZwf
4ZscqfNhNajLHzMAObhbYLpuJw4XjChAmwFMgoJqsYGxxntJNnMaQSV6S0ZqP+vyAqXIsb8BA7tR
dPZ0od25xo5FQuFAvbNMjHeYEurfA1lvPJshM19F1uQJTMW+YSvHbIPaaIqkCXgc92qpd4RVQaj8
l1BMkI98z2+3CzbdZHbCTn13tgkZnwO+nSJe+xET0GEUGmR8mBsYOijGMftt6VL62p6e40C0HFOm
219rAg1OcxvMpePASz+djUYLinQo2AbzAbkcwrbTYvJqt4ztpwmIqfoSrjcBRuzyVYgistgrSNGS
kkJKdY9mqOskPX2mcIVFG85k/xbdmvX7vGGVULhPVK+b6BSH+Upbw8wr7ryfatPwW9emKn92F1pS
q5CZcIR3g6RKmfT1BTTjEN33B0OJIbNEzewhOS1DOEUIdeby7DyZBchAbmRFEPTlsqbMsriyA0kX
qWX99J3A2NMbJit4Cipdds+He/uvEvXpG2WQTKEGazsVo7CFYMZuZ+lT5jmocSIfIs2s5HBLJE1a
WtJFzwNypNAU66bsYPphYXjjvYdb4y/fT9dfry8IW0JRw0uQllENm6+DtH4emuwsAboLjBSmLlS0
gQsxNBpsAHkwe6OyJaUZ1nTtNJDw/bwY3A0rbsn/Is9hjMBptYclwV/bhnhuBVZP8q1/30XVVuS5
tT0CS8TkWphhhTW8aFyR2e9L0o2T3HLHrGV6MEDr3Q9BYaBAf/FLdVcWGAmEh0P2hp4nkqtpqcca
mI/dTMJcpZ4ej1Tyqa9xV0btX2BCFvl6ENnNTzi6+esaoP97xt+GIrCuRkqw3BGMKX8UqXmzIBXx
XBrYJD53M9619pPAGQ0RSkqQtFH0DUTUh2S8mJTLM/x/G7DSqwrlqjwZ5OOGEIFmxpCfd24OM56j
qQ9+YNmAWYtng98HMC5xnvzp46b8uFbLnZNyAILu7RL39ni5fiHzj8M0JtQjLvwV4HBQ0ngyrrTh
gBCz83tTNKfKQI++CWsL+QqNRlgc8xQu/7pbzHhXF7R+v6mqB1B3Kb3DdOS/qGQESXTxM/fSo/vZ
AjeFrdnSIHAGdTajUY6PmsvcDmo9NWbpxjOe53aAZbxfGQxP54iuoePJEM8PBzS5hzgERlfy3yrd
yhQSunXpi+X/KjMa/6OkmlV1uGJ4KkhK3WOQ+FYaY/ds2weac4A470vQnYNAgSSwHKyQWQypNjJQ
jxPHrPcR98Zn3/YfiDYLxMkxDgk+BHyPRqjmgCOMU5DCLhtqkz7pSkcm/PGX0UxVfq5zYNlxBQM6
n/zFepr1kzegCH/aFStz2/6fDPj0sbazfXqSv67JjDxt3z53evYHOJBSti1N8hDnlklXOOME/jUT
HROzFhlMiCSBLXc9t3tv//snz3EKinTK08s7s9mmT/W7GW+zx6XxcCy2blqYaoHR92hqEYY4z4xt
chhtLEMD1kW7r7ZCw+eU9rTsaqcbv7ZX1vQW7KwxUGOzwl0ro9uTzZLmCjNzsbldFN6aNJccytGR
w2OuOarneKWEiN5em9iB4X6O27Ex/uewpQ3uWTN6Rff2s7nlAtvzpA4Nfd7aq9pRfI2C/NYI1DKA
DcahvOMeE5WMup2bhEEAXrccHB8VeDsqlX+UnOaKnpWti2UvuZ9aynCLRu9Y7r70bYRanTn4u3pz
aV7H40QI5xSkPeenCrUA1a1f7ceWxPI8oEiq7nWVYqHG2jLdyZfhVKqNoQyMOPP4KAGrcjgn51b6
FGzaVDKh1vYXgeFfBgsCGIIZxOltjbnLn2NUuniDIwho+krwLZ/jDMomc901Lv0a+LzOSAwhFxk4
zHfJB+RCy0EGaPuiYKBRQHKbXljlzxSq0RKc6NkcGBeGP7c0gF1xaQvy09+9In6aXVsgZ/3kEaPr
IKWDzi+Le53skpjmj16uMUriXLgtrKCfbwVhjxx7YmeOK21oZOFWMKNyUs8GrhAZRaHE40ZOriv4
6CRiH43N8uwB2u5n1SuqUe76/SeCABl/Qx+fD6iphRAhJet5FC2fKVYVSnupsJOqr6T8E5iOJZEV
7tnmZjsZFl+CeYLOobaLtUz+88ryLmx+FDygbPnw6C38Kq+Keg4aOvZBBhGEoNbtDfYighNQKjJN
8MeUSq9Uv3/uynv2gFSJnQVKehPRBMhsU3e47N5IeDdGBsS1vEe8/sMC8MOUO51nghXfWfh2/3FB
xlp/3lVstGsr0B3nA7Dth2GiaUJfB5Dc8NF04FyMV+WDOWDiSOLNUpNiTZs7YWwY/s7mo+JzL0RH
HDvyI1IQhz64jW0DTBZ0c9gMiyNhiCGQxJnrkduLZchOLXlZJLQfVCksDoqJ+WBseCXG+QhkuTtH
qPpju0owQQ/serrHF7EnISdAXs+M71fygcVqmRZbmaNbqczwQFxnmK648Bm8D+LWmk48Uc0ndP14
lf32eg3G0sejrLNUyqe1n9ys1CBAFjpebIUG4ppHeCsextKuKS9KsIPXUCLuw+ylEVknWpAx2POB
Y7HlgGJPt8O3iTFYBFgoZj0tQKtSl9OSSwX/JenDMtKQ0+p0SexznHzxI1Xd5T0tGFHDlI102Avh
ewYr8fQ1T4kmqCftj4yytDyqBPucFpKZZMpRxK2cZYZUxIScDhOh+y5sB1XcN49xIoD4HTfZ4VFH
PqIlt2vnZ3/A0zRaC/ojTJNAvfgMhcY1WztQXyfwcGmV5YOWkjm54tX+I0biWR2d1Db1hlevlMH8
ntDRYhZ5lzCdeKChieYnFlRQ7ZWNd0Bu5XY3tFKwmuyn5TOyLVHWQ1YI3dNsL2CXx51NuvKM+fxX
blSjcV3Jr4MMnUKgh0Qa7XqBUNDFTjtIjcIGbE93ar414QqkQrt2AV2j6LFOcb3/jVBJ0gXNq3A7
CVs/2ZnqgEdQtDPpUgOzRc6Wb62cWLguHcsWW4XmBepy0g8kPiZUo2elhPXf38ZJ8I5VS3HAGGF6
j2Fx1SvRaINJMhfG9kD6pWf7PiVf2Hz91Ei/W5FH/V9WX7HRIZh718PGm6KRcibhOHRRaC/ezkp7
wrraoYakUf2bhY+0938iMBNTLFuuzGucw+I7FVux2REjSD8QA5HWQOPIWzY1KEGLuv2U0opfaSi1
3z1SEL/TXQvDPCao/FdFml7uA03vUgQ46AddA8HOMrR0I6E0f9GQIZobtdbF3nBN+tJV/YWlGnVZ
tNq/iAj3e1yH7iAtszaIlopJGnoKy3X3gyZklw1hgsSsLXhXpt1hdycpalvPI1zm5cqvbXqCNE+/
HC16hTHChbrzfxf6sGscP4gsOxNlII0aIAkTQb7qzJg82MdFe5frToo09QU7TkU4WSYnAp667soA
fPUaNpXuT3b3Aq7nrswId6853nCloAwMuQkrfJz5ru8q3SflPTprfoCY+RHH5WNOSCn1djeiKyg7
bqiSJz1HNxQ4XZSeof0A7+T6QVw7engEkQt79nIYWqX1BaGrxak6964seXkM+wbAximhCzDYA7Ae
IAbgMlLfeAPoaIN4xsOXaeNRF/v1nFlm1UdNBRg8B/qaWH3m70UlBvmZDy6GD+ypsmyj+JyHjZMT
9SW2BY3Nm1Hcocu+UZSP+8UJsVgmF0Ypg59cexnOLZH/6XwnKoRDAAP2C8A0yIaKQLNigtTWRaeC
ytH+e24IXBvq+DCy+izfdxyYjWoZ3wMmhD02d8MSKpApA9Nli1yho47faLH0FIfIHAyrTgY+tY82
qBDCmYK3WXFFLZoVhUfC957b0MBHuZjJJr4B5lJIWL1aKdwQoAloSAdSnezYKejFe2pLhGLXG5Rx
v1u3ax7rVtQYBnjprEhB2A6xbDGEaBewIWsHdKip2Q/OBaODNsNe/4p740aPgEisaR6NlB+1ZUTN
WMrw+pCR5Q2Sie25qiQH9X2S8hdsD9nWPeqinRJrNWEvCSoFE78Zu36xvB0F68v5RsrVXBrHpgm3
QNtSkYUeQl8jsfkbYttg6ZXuNI/TTSvSuRcVUUM8LGl6sMY4gNsWW7kMLO8mE9nHDuXOpGSVt6Ov
374AwbJZlVOdRNue/RxCgV4FqP7UBws92IlV48DraPUhf5pHqOJq1cp6HH1oOrwYmLwD5kjXS8TQ
LI0zJUnTcXD5+Ni6ApqdlvXd1Vb1vdpJhXAwnZqVBenAqXXWB4Zs4VlMFNB1vQootm1HTk6GRRMC
IPjHTCzv5Hrz/FaA7n8BLJzgIFiXXYYU8IUs3pA7cjxvh9ZxWCwWaoRWl0YYiF1y41PMxW3mmeEp
+QG/5SOl32xBcrecj/MOiX5Sp1UQ9LiPVjXYzkHE9gdA3C57JIE14GcsTcRMqElZSFVIGnk6cP5J
yiNaXGKhmCxuQiqUwbhOJjlzrzM55ZT2jhLMHGIDWtUcU/bC63SGDbe/8ms4d/OopPc54PYs2ta0
6wFZocEiQlublx+qkrNt4E2mrOR2iy/hxyv/aue4sXVAjOROl12CY4eDc3f4o5p3deA5aRFFzkIY
fCAklKhHBktTOecXqQl5iaHDoTbTYaL2JXlyHFdg1y7cumQ/UJds2+zftYGUiCUNsEop1KezBoaT
vsAqiCKdF+4ozuF8hIuyahgR+m7XDq/FY3N5EWcrbAv4RAGk57sjbZrqC1TRU5mSeNwbXiFFu4T9
4ET+fP+9xxCAO/78+rnlPjw0LTQarNfhPSrAfgDiD+HqtjltIrxV6r5KdWT1Y7poQpZ/hFAG1YsB
QqCQ4DKNvWRMbs7jOQOyurBOCSkbyeKunkATT7p0xinjh5wgN5kLjIQeMHXrRds9lrh/k7lpx+PZ
uaLi9H3EZKOvxYPHv7faqgXEfo/3iQgfhf+Wr4Omf967mDb0QQckIiu06x34lJIk8lYgx2DzKQe4
y085VNY/rav19fHYtM4CNV0kjXsQbwREhEj9+rEic2oQwf7vkwFdbvf9ZvscYRJp1lCkdrz2B1gd
VGtzwo/rsovLfPjTikv5PNWYEsETgGxaU3bLdYOcfkGYBrr+G8diOCa+JMSxNSoO2O5t8qq1UgE4
2lFtG88eDdmQu0FSzgu2MgfR1IAnnfcDuMnnhyvNW7x1C8+sXw9uFTAMbOaJw5pga+fIYnCjQSN2
0y5IAJ2xtmpYSl7eafsEF3dejdO61iwHrOMn7JZt5gRPAVZWmiGOWNZmc2y2XZmEWBt5OAMHgVwy
ChNsVmXGwp6EpRMDSjrB+XcpzRrul9trXtrBFJPInaup7F2mNpddr1RP5HH2KIDSe3yCpsHaOW82
gjRKT4wShe1hawPV89SKFI06SfMkxkd8Ftb16jhERmmF+rRTdNQlii+mL2baT4SjYuoLBS3q+jkz
V7t8rvxKUhkLPLYTYiXByt2DJ2r9Ih0/RJp68RQEAzrNU6dzQ3JI/UIowATH2fDEDRclpuz6MXZ+
NsR4819E+pP0Y5Vx0XiG01XLr4cBS34Q1QI5g6KSozebXy+SdSOmVir08VI51p/mCuSAGz+5cnfB
2L+YcFYj5BZxSpiifko19CavwcK+sGoDgYfxJT1e2w0SGc6KeOVo5PJk7Qqk8Rs7r4KJGHx5GE0/
ilhzz9i28ANwQ9GnN5ldzonHDRLxrgTEp30Ia0q1DpDCAOhZhkqAGulLZ8C3OYH0NhBGX1rYcykh
bZQ9oepeLkB5yze/J+a7Dj5tatL9SnV6dfZewLRB5k8f0UeuBvEIFfeNc1ZQAnh3xfgM+Zxf7daw
xyW4VQ6zZCLD2HzAi6JupB9aHTrCvcFpYzds6L7ofhZMK8VY0kCLYe0s3B8PVgDfGzbiYe4XcRzs
XEL73+n3fvNAl4HNJdR84+CUiD9XksJnT/nLLA6pl7fLqbR/6MZYWNBe9YUBYhO9uNHwPYinRTGs
f0yi6vYye2wt10gvollgoVJphYR7gKWna1pfTmn+4TAD+aRTrlO8JEM1Ib+PwKaPYTE4WtfIOjTy
3g+8IcBw74aPfKHDwTwKRTRUgPH64zhxVFY79VavQYitRRlIGY8zlnpdDqdQw6gDuPgAP61djFFU
KX43KnUiTcXHjjVDcfse7cpTzDaExv27DH62IJWUBAQLAIV5PPK7lPqWV7lvIGLhPtkdsMjvpNiM
jFjuOEZ/7FlJbjxbmXhkGQPpBGjUqNAw6xi7VJkkZBu+W0m0aN53P9eVlwqra+H5cza3H3lyog7x
jke7Dk4XpVX+Ex/4L/lhcDoWT7bV7rsDqcsNSLkb9xF5gmdFHZp9oRGvbM6KvpJLVpgY7h8S8MUP
Ty4mfqJ19kAKzQtQwwTuQ7rXe8g1PYqhU52culT0NUCJ3SjcbfKyIyY+RIDmN0c2/WICC8qiwS2t
wu/+jxXCM/ShEnRMa7AxmFojPH3sHMe6ESlCcfZP1+mknRqMJVVqjUgwMe0BJd3OQP11wSVGYfpo
OR+KCTNjWDE9e5ZKlGiZkwFHDUS+zso7ZW1jW2kiTwO2uIUP9LLStY3nlkyzlJ3LFQukREeZSCFt
8Td17u3vbUfFeo1eHv6Evy4949pvOK21a25nv2KhHusAyydDNTMr0aVPHEuigmEYwjcAWJGUKL9+
vRwo0BwuabL4Vy0XSikZu1JVeaKiOzF8YJsDCOvfstFUC+lWWc+zSjuaTQkvXEBm/12gXNL1gFZP
ackBVyvYu5KRE/6KrDbTy5AiLL41zUKBx05K9srEW7ZwF36KVlpBfQj1KrQGTGDq7N/FS2Heet5J
PGMC813W78Cctxxc/JUgNCHUuBr1ucjgGzg37gNqcAsieBHiI8xkr6pSn3qWkQ91C/zwIAtkLw0u
amE9c/KNM55f9dCURW8FYuACuIdsXpSOCFGxA6BbeFvwIuu+M/tF6FLJCZDekd1h40cMRyuZhALf
KCiJCxBF/yPKn3/Xbi+dUbkbGhn3X96mSgkxOuAlhTf9eDK9r6QmV8sEYYN9dUFT6k7vZ98XhPAs
fQSlOh0F6cuMq5+k7vp7ajDS7GrJiaudRyze+GV46vLJGVpXd9yKcB/hsLHrGMbWsDDsSZJuyvTy
QiZMEnFg2Os3dyMPZl58Gd4dH8xQx0/rC7E7BFrX9qVdP9ia9d/ySViMVPC8lWZ59t7EccIBdHXz
w5wQTi03T7dun7dbJ/Unzt1/A6eQUlkxjZX7/AB1ySeV4Cr22fu4JcDcH3BGbZeOj/8MMB7REK2F
SGrmrg53/y9dAEcCExVqIMt3mfmsblEUJ1zKTmSGPsklYOjbl860rp+nnkoHmwIUWdD9fXOFvcCV
KpzsxgW4I98CiG6s0gaqsciN4hFh88VTUyPmaYf5oxrvkY4CU9Rsi4X6t356Cpm/fxHHG18lgOsS
gZXg+Km5WaDkdy1S6jB4Ch36QoAUIzoby2UbRSPJf652u3sUP1QvyUodlbbN/9+JtUMwznIo5f8A
k2G2dyMxiYDPI8ocLyJhabnkiWSvSJFAdK4IKMKB4OpaTqE+fixqENN9xal/fsD56sAIIiYwg395
0Yd9cBEDHZU3R3A6cE5H0NTllJn80WlACGifaGVBh2opTqFvq2wIsMa9ANsjnMTCNqZI1qyHkxkg
SX5w5x0jzx/cLoDab5j2ofLWWZwbkmT7ppLgSorlGJYx5K/Pmprg/gM2Zetvw5bUwvC2lXzZfp02
T4nt8yL9sHsW3949yDbBIoIRxbTEDLKrpX0O22pmLRWsUJ65DRgNWZgmUShsaWXT0GJeVc1jWki3
rpiUzwnWzwqkyQPvL+uqJjewCvEF6gEAHt3zeD2GNiBQAFygGssUrJIuhWI1pvW+tarsCRxJSGvB
fszkeGyEVyR1Klt2+Do+3mnnvUw3FiFxESP33NAvbTrHV/0WwrKOYkEwMilAF9mi1DxaaQilT3lp
7zO9qvzfEy8wJNMM480/osJrQrWP344vUjQVY876lXHPj5AH4ARTO0NcG+jyq8HfUMkhlSSClGno
9PmtrpNCh98F/mWoTChakblMEkWyfe5SBct3bLxnjx9L3vLXMhXWZaIa9N+uaulOoUuUYeCmWkzz
7WRQR40UKFZr6dBpDyN0JKS6cbQ2QvWH1BNuxcMmeAKva7/+JPoMOpMiOJN38O9AEvfr6/H0YcEs
slUOUsNKLrd/hHfAs/vdp0cXYPikggFQxVihtWZmr+0UpP4qQmasd9ce0X5U7VaE7BGStZVGFRSq
jeIbnrcHowCW4anOF6Nz5BU19ILnNvzoDQtSkv8Ck6tk1b9bhvKM2eUWQEzeY2qX3dSL6J6OXuRM
dThZ2PK9Dx+3x+2gtDZ37sKJ8kPOL3XXV/XtC9QpHRjEkmVEwZqzX9Wgo/WJUV7mCqedSslw1rAb
Tbk2GVAWLU1BfUPUd2ViJCUKegu08jUVEdEtd2tjp3rC0d2TFd93rqIw4h2GuQlybHScZzwpngPy
bTjdOe/72vk+5VSgf72SeYHGyNORNryhlHhGdp+CNcQE8wRhusFjvGoKV4D+PN1WWK1RYJKxLPdD
ThK0m6z1zuLFew5W9TmQwEG5m5vqv76fTSHwbfGkMSQtR6wHkleHiBWAKhKkAq3KBuH0tySEvOQb
eTBm8zhwIbzfDDCEUCBiniQfmkVgAcfnp2VxQVwr0vhqqKuxnzhu1Xq2FhdsXdrNHwtzMvmHoqkN
fas9v5x3FZzdW3beHqZ8O6Ume86HRdYdlODkAoYTHLAbqUwXlP6k2CkD4hK7BCGvGAFdxBzzsFYY
rIxAhX1XOArGCq67XUfgz5TsPA4W0RNapcVmMP09DxSd175IQbcNRPc5vsKvpt2IrCzfEYhzOAop
6+pw9DWDal8zjIAVVo8yK1hdtOOh8f1Gq5XwHSYE5jtbqaVAO8YjYekwwMwkD72OFxsazR0eVqgT
+7Dm/RNYzuV5Z5yFIB3jHh+WEY28YL8hVk0qBwY1OxspT8Zt8AcywEsMYi2JxDvRbWknbwKUucC0
03x9CadjkdGw4R1yjrha9e7ppTEdeBurO5aLO566YlAoUPtCdoc7zUpkf7ihLwuJm4Ru+OBwRI+/
tC0XG3kahYIRANhXXGkLdFdWQJpEpaKh0oyWcmZEtsraAkt0/3zkAiyIc9uvPJoT3Q5opzCj2azm
QtpauZ3xYFASaPbnWT3YF1DM3u/7EOpM9XR9LxrceJi2yF5UT9JndgmOeFlOjSGJed2m09SHrBSn
51H714hWOmFXZKkQgLevjBf79hJ8kCO9GuAf5A5XF78U5oreJGdnJ6KSL+jAR2X7UzOp4fQTjhlu
srsuAe+lcbeAy4dnCxt2OVxAQXgKMWno0PMEBz1QY2pTCQGPC/EnLz9i46NO8iXdASdsgF8C4PLt
eT0hr8pkGh6jaZ3byvdm6hjuqHKLXJ/8z2cE84Pbj+pK9eJBVlXankOolM45dqVjiYGiOgaTYXQB
PBNO8g33vd2vXI5w50apOV/lnUyZdtkOvASKdwIv9D6A+zVI1Dc6C4FsC/miZ5/DHcflAKDxgBAe
o7gwLNQCVoL50Pxztg8DNeaV3UmH6QkJvILbxxeE7ICKU0eESG1pClOAEtqR/yG3PMFOWbfMmtul
u21rKk9tAFXAe3q47Ix//9aoZ1zKF8mBCJlYoYSnXC9fr4MIA8VvrbYai5ZKyNvfP6qiPQefwyL2
ZOItiWOMQ5k2YVqY0VS3K/bwmRjwmDzyfcZBe9uu5EdBX0pu8E9+V8AGS4oqrLJGUwvnSKOKp6Rh
LVSTjm3icShLbnSl1GoUuR3BxGgpERBItPtZIbsZFf98Z7/URK6ZkeliLuxFgHC9re8aGmKR4JEq
zBj/wj69QroeJbLK6Iv166uR6ZNhE6dBzDG0FCSZ0iaN0rX0+MZGfs/5nwwz9Uhq+cofZmPDhA1k
/px+dCY4isgDAN7ERWmE6+YaHi7GP0Yq/TNZXTY/KFb7YCDYL7ou8oT7vS9KXVzqONw3e4K0xxc9
O9wJzzZswto4OuiusX8q72bVC/Zyp9cahULtJEM2udCp3MfBGEyq+O/k9OvEPo2nq0665y53RJY7
wa1elQKjqmXCqzpgCgJskhXYEUWVG+zIXFZKr0qirkQpZTuUdGd4ggc4KV1nGo3+xgJ1aHsTBr8G
k7pZsKoY5OECEahcQDKX8t1koKGVYzd6MLJvvJ/Y1rFnYiAoh85dQOItRY31fpSv3YMtTW9/ROTM
EDpLRT40YosXrA2IJO+jARMSIm0Mk+pcOCCkoGtUYWE7rqDPwEw8dGNcOuCtx+xvvWVKJLVLIbqT
mGmcJ20uAeTv5o5Ws7YWlJRAAC1HeMxIE6msZDh9abK75tqrBN6NeoQE663QdThZFi78pxYYLeTu
Q6nGZCHdUmc4hTI06+8u12IS4HOE6wMRFdQfkL0f0oADQ9jgU3LzOL4vFhKNiFR1YzwuEaeLDvio
KFEHd+5KGdxZfoANEg9uBStIl/vK2czWHgJHBfiOaheQgCkcAQT0j4IncgvYBdq6Zg+Amo7Owdd+
ZFhdNFJUp6jbpZG690TgCLdHJFQIOpwgfRWxItjl6WbT7g6yMrm/p2EtayS9iXpqcapYnHd2v+9J
mAAe1PuONLWrC27BmCsBNJUjfML9dAAbvjDgI8A50xzbFVvyxeJ2F49/Ezdlrja8v/7jkFomPejX
1qfkgv/+gOzKIvsFLxktVmXY+wWitxAyMeeZ/8N/3ixChR5rdn4q8O1dt63K3P9k6I20rqja4ZHZ
eeYNl53Xvnr1lcTIY5HBJcgOueIOErM9b6FL3vkIFT0t5pVnjVKS5q8iN4c1/wYIOD1HRJUuvXzM
EW+Pm+lEnsF//BW1yG02SHMVvfRjn0EBIQFM2ABPVx42UdgafSQS4juQgwXESTlEaJMatWVkvtG2
mguMpoaPXji8PuIhZU138pVuwOKqF4ZshN1VlZVjigY6OZxaoRIwNFNSdEtnr/m3agoPr0pWJCUg
JZxpKTTrdH+tC97X6H3UjAYVJOV9+YNrmV1V2fJtulHmIHKrVzsCdoryGiruayo013h08uLrVha/
UCQRPQ7jDZvEoiw5FGZ3E/gaZIFR4axBSkAORdkC1Aw7+cb92rM2UEbc6tMUzDz2YLpmq5rcJ8Ei
C9wmJZ/oLN+PefwY3Fqi2V55SrpHZdphBJo+GmbJNzDzvd8RSLd9d/73SQVUsURXFAqb6MfvCqWs
6yLAC0NK1vkZAEx8sFbW0EdMqKf+zVe2YeYL/0JPSSYkCXneoJYe+AH+pTw2m0vDVxWVoakHmmwr
2qjgdgbyCj2aruBzUt5O5zCqSLyJGj4yvFWH76pl44HP6Xy9NbhCwywj2SfroF+TeMcYu0xrOEzU
YJwlWm8w+GB277Vxa7Q/PjYXwvGHAUKbkNGbvfysASV92+4evSrja+AgsU7D2rbKbvZ+btzUyzKk
7vBEEoMm1Y0maUXToc6LlJCDcsXXwjlNzvDPTjrXpb/yfFvsYODVWmfgbZLSkQ3Y42wbWiQvyAT1
Fq+IuS5x1ZWOU4/Vq3pwG3AwSrLNka5uAtfLbWDTM/IYDZp2euZclzX2yrEp1T+SROgZRW952G2S
Mgd2dji0dF1KX1r3auyvzzOfWWfCfeC2ev5Iky+h1DbduJniKvEvKSrcrRqX7vj1utkQxJCK1RbT
bVRm57KAOLFiL/SGZtQ6ocMuPT3Pjrk1aWU+Ewu8LpHasKVAFYfit+p9jkw5cdKRxu2JH6wTK7Fg
MoSuHBjRtp+eM3MVqfiu9aKbKoXcI7Jaexe5cykCqF31/Z+OsIEXjlYpydTHgoHjZ51nh/q8t0o+
5IDSvhMGk0/paWSaxMPWeIMNmTM5zyLexEgf8Q7FPa5dkjba8B7ijs8jNPifzpM6QxmDUnT4181w
IMp2jV4Qsm8RDNVEpE3ZBArrLV43KI62c0nMcDlAwukJA7JO/H/2d+Z8h4FuXv63FyuSXsWPy5EH
HHkzGoc1eIbZ9IEUy1XdWZ4YdeGsdmEG39He3hbG59bplRGwP3l8gGAcSun2j64F3rY+eJ6Qz1Kr
9hAeihOWTfjDbFXX0+tMZZCKADGh8F21JR1obUt1mgpeF5rdvlccNAOdBVN3ffBJOT5eB4y7QIYs
LsO59SHWyb4iWS9xbzQKBIjSlwj67KIvlb4wF8dBFJrHWrT2bVFu5AG9rhvkF2Xs+yxikP8S9EES
w6gNl7EJaMeW/aC+Hye0FlCjG77qkNS5ZN39SIw5ZgIiAJX+4zzDqjTY/O54ulEzV6P7k9r06VOy
QktZknVa13M97cXkGZ7ed5XseV5ucETZ3RPTS1hYBs07h9GUpZsPjC+ucIsT3NIQjBgnww0VelsU
hbg0RP7ZykuOu4q+qPwV2V4wnCmphSSdP9BwPXmCCqEz/hzqqbMAwzMH1vuk1cU7Y/t/Xz/bhXex
Wr2Ij7DANEmSRGHcp7k1n4Cnsw//8eaeIfh5NjotjxWgY629rflzLGaV8R5HvbJhdPxaMv23SsmM
x04eDXEjY1gQGFp1KTBJxzUpkkVsPHNDgLSlPI1C1ljXcxn03riEaQ0XErnxG7o4x2vvTfhSh+s2
5GmyLOm4iRjfyC5gvvVEs2x9UPmuSB/3z0YFT1Q4K0m8xd0ZX7F6jLlwOjQe0mc9yWdcanyGURqR
bZhZXHHukDJbKxJ+eCxb45naQ6WW7UJ0XRIzPlf7+E2lddeeNp1eTBPqfiPiqrMn5Km2p6l5yslN
ei7YlG7oSWIisaH78Gzf7jirFTdXdn9yhMf92yY/ZFqPQKPFU9ypr00mRVQVQHkJzEaDo3P7pbw/
0SHR7eQm6dfiNTeJHVzLluE0IeKk1LS21dhPGjgz8SX1NsejqKwwlOHURAcCCCbiC3li9Fo4AxjQ
u3dnjOvegfbkEKN+3wLIrGxY1Eh8YTII8RIo4ulNj9NxIA4nX1JL3e42fj6SlG7ydphxfHpLdY5l
6YzyOgfw+2KAofMsXrHvXT7bsrSk8atwleEprACW6OwLp/NuFYfDlB76szvbunVXp+Ub97qSwLLB
e8jSxovoJm10ge7K3wLOwgOQKzx8+EeEECNRBCmUM0h+zJm0cznng8oYYMnft4DdGj3HS33GZUjj
43xhoxQ/hMrq6OG/ip335wuNvMbN3iOXBqorSFpPvuUG+aVmv8QapeznS+AYUhtLpfsbkWSTBH2I
orNaJtWy6VpqDohnhIIjwWPoLqwbDf4zPIj39KqHlOg6eiig91soVFISa/b6M2HVsUoDufHVyfjp
eKxt6HoOVQcuTvrdbWiX1El6eh9C/Iefw4v5rfzrPUZ6vIhiSzk5ITE2/eaw7zcFXz5IX+DANufC
TF6/jCgZc5aHjxsng3RgaoHbJx7jri6xusIPa/5IZyKlMGqZXp07HyOzKC4ntnTMKmTloWZfi4o7
0ypvTRC9jZpHcFKvqm6ySHjxjOq71NmgvfQrfjqBIUGAOPPWLsh1I2FFnScPN/waZrYBBp90XUkz
4RkUyoQ+fSs4opzoTjOvdVsB3S+vTpqEEDRYa53Qb1kmmXTzANhIcxni290LCk8WbXepsjE8MqLi
CNge3dpNIe6aUiEZBZVsELDhrwnTdHGb2WkRcirvjpjFcQXOGj4ANyk4oTXhLev0tEK+BIxrZcpb
RZQytsh/3LZKdwkgXzG45Ic1uX0D+eTopoamnAQj3d+B38Dbl0IVdT2MKY25ig78v1klXfkHVJUf
Kr6g2WATL6t46PKYF4j1hPQTnKQR1OYRRO/5VtWUxoxUDfeu1/k0xxyVhv2IT7Joa4NeoyzOJ6IU
POzpik8WVa0UJNO2CBCEiLeNMx6AN28BEFY735/wFC9FjEgMX2mvC94ZHHh3j2A0s7RoKMMjTZWG
jTKrtVQHC4lcxHVk4zLkWHTWgT/VaBYuBqiRHq/+kTk5hBjxLJIESU2GxxFFgwi5V7EZroFgId0n
81JVcZ4syN07m3fi+B0d4DfjrOB4AmA2nO5aXTRGpZWiZYLUuKxbGVVvdamoSIC3y5G8V3qt1vkK
my/H9T2TNDQ7SVeP3zcttC+Yl4rG2VtFLxWfk/qJAdolCOQvkTkc3a3CpNUFUeU5i9CPmW+fFeOg
iwXqGVpgCxvdiBthiS4yluIANgygIEtyJuhul7sHafeKoUIv+UUzTM5gfmiV8ojCgmjorAvZILkH
pGofHLIBdetrnvI9kk4ImMaQVPI2NspF2hrjjamfkPtsVwM1xxjtop9ssaeiCOESwCD0ZIo/thrF
ZK5yhmp5CbSVoAvnInFzxVwfadVNyrQs46/DYM41XdXQSf9I/SsMbN8Xe91ZW3qhOclmRLBH9f0e
wSmWs/uyGA4NOVg3/2C0z4ZlyB06bp1TL2ab2H+oLx9ef1ANW2iXsAi7ySmqMW9g2RpI7XLwNy9i
tFRFt3gzv1rJm/Un+WOjEsurptR6OwWlnLC7eDhCazpAzuOXE+t9UFdbXPKgOIRVu503ACT83CXk
AghHHRR2VvMQClBwK9FcGbaD9IsPut+EiVhTHiQsWm79QpRO/34Oa+k0ffuQT/TQSTSIy+cGJr/5
l3dhp9LU2E1iXQkANcdzGvnTjUyq8wRVfLFw5kUx45AzUYYVcRrSvOPLvewI7WoMxklj95J5tau6
miNjfVNTiYnY3Us4ElIwDcBJ7mALbvNrT3oXL6zix+SS/X38AqkH6gYa5Qa6KDLabKV7UPpCtFyL
2iTBV8V9a/+GS0Yp/VLDhmS491HOLZu2+5M3zYk/vc72MG3W9Hq65Gul1Cj/rWwIku4oCHJu6NTY
30cdTZTUv5qBNRBCUV7HdDCh+IT5NEjLfqMG6+6L5qiPbxUV4cb4SlAnlKfoQvXSvbbHVMsIrKe6
kmtpG2QfBdOz8zEOzJlCBQg5TdZgwyJpGTjPf8Xt7Del0kGrhQSQ2CISk6u+GOs68VV3WIMQXvcf
2S48fyBCI7rG8jNx0oRJ7aLa60JcXvVYYuM0KsRt6qs3fsA0QMpIoIVgzRZJT6ohdfCKqhQ5+diJ
gSXE09rdvbFHAVurGbbDVm25nJsaEAoCm96WLNTvGT0tOJVUCMWhWnnEmX8Yd9qd/RAABlgprSMe
rCu1LG9Cgog9xclQcef6+UaBadCuFZlft0NvnMRYsg4d7lvhSGEmwEs9ec3HK5fUwAeE1jsOcjcH
PCdWWxgIXOl9tO/yruZzmitKRkjFccEc/7okZuYxcQ0ul2sUo/D72z+r/fIPmrt+A+YqbUcISLp3
D0p/LwH/bsZEYVuwF6vnxB2Kiv7+RkLkYSORGjeZ8uDDaobKDBy0QMibLVj1QxN/YxZkyhUZ48cb
FXOv3mJv5WMt4m3qDkrqSxTZqoXtkID5ju3GQ33X5TE9MhDZcxPhlx/DpNFLjCdR1BB0m0Rb319y
DLc5kDRBBsKoWbesSWu2qNoDqjRoI4uIgzV00IOOt8Y5bYYRJsMQl0UHQBb3phsK/AW5j9iBJbr8
vcBFtIF2BWKIMkKD45UO7Q6rtKenzyG2wxC2C30LEIECHBADrmJ/db0t5Ia2jOy3fzwbHu9ZJDGu
rPBhI4+RrGa2advqSM/dACmxjnM5VNEg98rX1afheHscoWaN4uEVdGDogN0aCaWSBhp9DKS9BHFw
Rur9ZtTsHglVGeKlgoYMqjOgqD46zDL1CFBjPpwNmv7Gq8ArrwtLew+UbcEJ2srj2vXtSu9odmZJ
dZYXG7A0b5At84bK+wTtKxhxs7eCYoyOG3HVB7VD0kpcVh6Bfh4GMwLrmabJIVggSQMio+f1Tklw
Z7BJAW+qed4su4Wxh4z7GvugG9N1M2YOaysZyjOdgqRN9538JEZejiWRJSD3ySwdmEoab/Ea8gFn
d0bi0nPRdv1h2S+OR1MFdcjEsKlvQVFc3kLvUtOcGEw3LC7cB9lGR9wYbbYVLPjxfnS/3wMxx1W2
zlAtz3MpPskxsCXcOWLb/7kkjz3TjAKzstN0PNDmLaYbg2ertv+8n9GxHrPrn15Sc21/UlU3OVF7
yKdTWRz9mIErLLA7qk1C72fOYIT5jGiRbTJHGOpP0e1qndHvdl+RAlBaRX3j6eGzAxgtVw3Eljtp
zT+C7ptRQH/53JIElBYicSh5aFCxj3w1Cpz7n9/DIRk7a6pnXkKRn4ZZRnqtY8gTHR4Kw6o3rk3F
C1Eorr+87xsvSUSILCBo7SVIsalgsrRvZ5470tWTHONNbYHRSUEYgKRCarvueMpVPevPasys+VSh
PBucM9dHUgebDxIhFnuuuPzdUPcD2O0whe9Wl7LoMK2Upm5mShb9W/YuyMBTY6j4Itb+HtqYxvxY
cX4MsA7YBJnLlIU4FTToy//iHOZfrDmgSpGUzCUIWWPnntAo4Mem0HFfhw8B4uSBqGTekz2LIY4/
hsHqNlaizcKeVUACpS3bhEzeIbsHJ+NrkaP/SBmVRB7LZNVGCrQMscDIHRNRKhatj7ai+9JVJob6
Wnnd8e57yDHjBCppDXCcxg8RgKjtB713DljRb23yhiFqcCtzHI8qvFmHg/ewhKc6SNtzFpurRsBv
sxl48oP+ADigVF4nwbTlW5SMVV9Ebs+vzyz7WCgGru7JOrgYdX8smIJrudW271SrK3Y2uYlvpgyY
5R+VJCGDgrZHT8XVKV/s5qnrylv6b2+NWGIF0TpgiRF8RC/vTEBI/JHP5pOLmN6AFt0Fjo6wnRdF
xyRhtxVBNDOPathewIU+MXjetBVMDVvXEub5Bbts8POBaCCfXz8kExLVwFL3/GwyjkPnZtj7S6kU
6PTEzMn0SDU6q9mTYqOHrCG/hQxGwdJGReclRs+z/RpMosgAmK3jWxEGtlTXLbG0S0Zo0t6yqXLL
mcUjpicN2jQADUo4AU8oShzmWsMW8rlUxjZwobUMXapv0fO++0IErXGnOfudLbqsnVI46k2bUcrd
A9mhSVzk0vwvTsPu4NwroqHRg5B+E2zjnVYSa3qv+kaINUYh5aZkbhSvhfPWL18gBdrdwHHuyQAg
qppuQpFliesDdz+Mx7MgondLI5aVzo0bT5I5MPqq6EqA+hnjjN3YcrBcuqDVRvZjZtGmp7Yt4iEo
hJFNGk2jr91kb6SDPBwk+HolvDYYgUZ0qO2i9k32Zj+0D7g0lTnVL5NbzklkyPaBB1dR3W51ZUoh
5hCvaPpF2fgc7KUwmZZ6YZSRUcrXvNNngB1bgKvPZyvgrlvl7afmW3oIeNarAElatMCZFgN1hKqm
dZ3rFwrB3D2SNIvgQgRrTmW7SdySgsUyvo/lm6EmZ+xQjSlKOCGkwRiFpp51O1xatdEp+zTwVqPk
OnymwI4X91raT2t9JpEWaLmPXx97Dzb2VvbsLkcdzO8gcI2Wfg2s+65zWaryUGgduc4kKFW8KZMG
JifTtFsP/yUNrFH9IcrUM89TO7msfYfG6gRqBs6dWJl0P49G1RpRN5CU2pfxtU4aQmEBomG7QWeW
VHzE4Z0/gu8i9IXtj3/629Nia0jcB29U8v0q5FVz6ffxcsAZAHMiGWluOcCTAZal681xHWVt5IAb
0PzoK94zAAAyhjlyAgBJKtUBTkVrmBTuuuVRectgZ83ZxL6v+xBiEKis64lCsXiIYugpcusD4MUT
wiz6AhPhztLaXoepf8Z8G8v1GheOlgzE+OZHvdLn1nGB/YsKwhUWT+7rlJ2T2JoIAmq+WU5TVIUw
EzrW6kj5ARz78kjz+7+4DFBU029ipQdFqwH2tTJoWqv7S715ZX4XffznvgY63aL3pT24vH/L/qJJ
hMWvRvf5C2ZQYCBW+0rfWMhGgEkFzZDR3i/qu+wRP49izBLplsf8nIn9FPW4hw0Ri6QRaRWDrmsS
sEsT8Al9AejiuNL/yY0g0K3FDQL91S2/el9L+DHulTdCVJvy5qi9zibguKIMVMGyNr0xAG0LxcaA
F0zvLLGMDVe5JU7at2KY2s6jagWFb1cqx2YnNmaWuXKmscgS7VejrhZQcEVjH5v+StZQNcYV7YQ3
chlDFfGP2T2OXhyZr28GpRlupb1jKFDH099ayktY8xXEoLUYljdnOmtTLGdzgIu+ZSl5/NU8FMaH
WB1Z7wlanLI8rQL/gAZTgB06zA97GRg+cGwV0tEqBdwcBdHiCyttQ6xfthh8oB8/MqYHK9h5zx12
XQXsxxyZSCAkkfVLFo3bxVJ4JLkQ0k/WdPp5bE/NKe0tRHwdzYegJU8Ha6VXTMyD6isclrXK4R/w
7bjMizSY3YYd3hN3K6pZ5wNl6JPMExgX7MAn506DhGdFBPNAv0ILqG5X/Uqvx+8o6yDqW+O7bsOg
vjY3+7NAmm5Z1gWlv2D0WBQgMZKbKRMVJXtb0bQe4Kavvsb+HkTPetLf6BDCMr9PHciG6BTjhP96
VrewqHxWFYHhtzIWDfNYiAzRqPdb+kjL/08zkpOaiaMoPXH1dpIKxyh0iv+lq1AyyIMhy6DEc92g
m8IsuiHqcxyn0rTH61Hw0s0xIflAzNpC1ID27sViRxxvMCOAvrPu08CWUMGcF2OhhD0NcuE70A55
3XJDSM28eYkxuB4R7HJglUQn3JBl+T26mkeKaKbcAeFKGJ08qTPjZ5lYZCSCDi5oanlK5zktauou
3jZK8t39+Wr/Fb0kOPF3go/8PdnZlzpB0gatLkEkcq3G02TA947dY9U4loC1vT/cSSnIt073bvNI
yeTOrz0vteMB4ddK9AfOFKj3+z3vW8FOUujuSPQMvDMXwoWchjkBk0LJCapItywP5YPUKFGuVh+r
4ZHpEEc3uMelNeW/uie+2Ua/LCBEHjd28t9USzJe12o8a8QNbSmaBemEv4V8yUvDYqRI+TjkdBtW
fEV59Imcw1h+VF01w0FCwN1ydFc5MNU1mohA4ZNarnXc7npGFWOJdjJAZHuTPX8Lh1gx5rKFOix4
uVNLhmQX+fjRfhYbPDB2DpYoZ880lEoTedLrFZupI3VoKy5AzxSEU1Ti6ykYfjg3IHsTtx9z481k
wRpkUUFi1RBl4ic4KcsW+Ofl2GcQ0ik1R6sGV0yzOAQvKQpn/ntFumrgfJJXotGUGOrd6VQwlz1V
8/tGOMlwWPB3bXRSrBHSG3TkPVWE/2Dz78JEm/cJAihuPAhOzKi+uN2tEJZTdv4f2wl5Y1ZnINBl
HTMlmrlLykAwLTPvWfPQpy91crrTJltv/3/+gCEOKmNGlX/rd3dqNLxnMpdYeRqBzXlrML06MsJB
QFrIkFKhenQlyrqIjW2ithJ0jHlWOn/rEbmqy9LJdlGjxFk8tZfuEEwiGd6TkyPWvop4BxVfUuCI
mS6cYkum9Fmr76y+P7t5N71R38w+0NUaXeQOGQg2xONvilyiyxiFv/lbNiMHkk5oIvEacpFQwxDF
i54f5KQVEzHuFG6QnAOOlGfD9gEi6RnDbG6Vi6auX0EOPgFpWJNcaAfOMIZx/YY0nfS5oEeNUnQX
YPJvZQpGf7fgWpGONOX9q1BhWNXxwPIuoqG/kdxyiDIn5J6TubSea8IYZynxht+6CZAIy9N3z8Do
G9Jou3I5kImPatOe667LsBniGnDrs0Wjj3KJk0KHAP1W42CgTF0UfnnskTmnCtptYp1IsZIljiRV
na505KXYcMkArucFEdP5hsUAs0511JCi8fKkGK7zgq24XbGTqy+3CmAnshmNZwh3K6zygC+hDOfM
B05s5KQZduz9DYzx5Yv2C9wYCE7QWJPL6Ux8uTm4X2Q1+Ovs3F0RFUI4rWhM0RwfR9guW3YQ0O1O
ypaJDwzRNAsCriegRB9lMhvtMSJNtvRsmJ2XycEd8HRX8c2+GaxIi/YALGwLan+qisPP+EQ5QMGa
ttuATQ4kIrM0nlVnZbuyN2uwM1+EmSsWMUzyatmwdA+DO4vusDmork2X5TTx5njfMV+b7zuND10C
mgVM/XZ/OWHchTNd44D/pa3jsMUPRCFjTYFE6iXigGbA8znD60XiZQWDi19Z00KJtx+kghzaJ5zu
Vx4E7sQXuO/S8DJwFtPyU+Riw+VeRaORiq+tW/tcDh7pcHR3QG00NtRHr31ACcleHYaXFrJIL+JH
mCgzfFS1jWTbPDrozmbrxSAajIU5SW52Dum5uMSqGLwYuZT8tQM7DN1P/1B/qNQNJikcoqhR5Y39
ZCtL7G1RWhz3+4dBdDzyxaRpvOVjU/+E/+VNcvaIFRZPfaENIzgPLJCaKrTarxfzWOJb50aDRoFa
5Gr8P1Mz+Gcr+eZAeJuQJaioRmQCVyyP5yfgWcTdmTfLzCIxrKmjYcqQXrGvw4zS/uO6xETpFvuk
Mhu/2pkqk81pKuBj9NRAevI7TT6FdYwcQXkFX84y9sLWc91oUQFtzij4RqBO5fUeWpbXApNcI7K8
6jWcRKohFgEXtBlifKkRE6gMl5RlBPNztag09a3vNYJOgyrAyyeJr1vNruvQt5IlGe9+wfnMIgbs
V31nnZf5F4GBS1vm2sfxa2h5UWS0Fz3BODsIwCcU6LzXEQHvYalO18bgqFsrQ8B/f4pA9b8rq76s
ClWWxuQiakICxIgpEJI0mWSFWZMnw3yAa9nFJVSm/fc82YU/b2FolEhz8/jjzF39xTCdDmcPgSax
NttAkFvZVWJ+oJ7eeNs7wbvTCUFuw43KExrHMKqP/bwoeUK87xwgCxQAzB4NIvcKy4S8pI2Ks91X
ztcl1Su1oMQnk5os88pRoiCsUvIXwj1KI3pHW19gMBAqtiSm46F/qfKY0rhodExgT2nSEWho9wd9
RczdATPWz/PsRnJRQXaUB2IRdFgF9pmROmbFgTeqblvj8NVwPZtIA2TKauIP59x+tFxeeYWuHjYT
t2FqN4gicBonr3nNJGJVsgevy7iadVqQSK0Q8OIIcZ9zfsLFNAasI+HMzZJcxuBZILk1dnyKnO/d
PAUiu7EAE2WZsCFNWkH0wZkl5T7B4yqfc8LvNmN9cAPhFiAiIeUZ2mAV6g4IIuSKLJ3MArFqWATP
hCLHnjkdL+uKFeQHEES074x7Sd3C1TkQv6nOS28vQ0m9ppd7RGgs15cOmpOT5mfieMXyv2ORCtby
0xzJbBDURs2BwAfbtWyeYHgrDkthJ4HlT3kV/duFPLWA8PsJXrOZlqHtclwzRUn3HOALvfItd3zr
Q++n7G8bzRaI/llMFh4MscDmW8cAYZu4ZModZPfCUaO9YycFTrquVD4aIQwMP0l0mffJaariGe8a
v9LqmmsVS3zVUHNEYSF4xCJv5W6xyIfADp74LRfV2+0Ax2URFOJlcZ5UN0m39Gza/NaLkGxiyOt8
Gf2/DgzyQPjc6RIJznMmaSuwiia6U2J8Ij5Y9wJ78pt3c/6glpcu/cdNztnKdIaqVsg09zgQ0Bo9
qFF0TEoJJdxYJR/rJkwR2Banh5qs0DIA9IiQCjAZ+bGT4O20NUmpMlyKKaIVDMnFh6mX79vYYVj+
sY3ofm4AiQcMuuY5NcGD42+c1pWdttM5pJ/Eq1dZNTo0cZK9VqZ2mcx7Dj65EEVOEO9m6NOPJelj
44kymJZUDWmRyFc1wIhQTMHmBGNmNgtPTVMvX9aUw3EEMslZME4w8opHa9Z17JBwlT+MVhS7tgLL
7hSylg6i8NNYZCRdRl6DHpH62bMU1nOcTzyhghpKNGh5PDdzT6FEhL7dhlDzUtI5L7r8HuJNFXPL
K4GrFQzOzm/6VSupVhWGjzdfyA8x8QGTC5BOKwm8/9iKR6jn11hR3vgzneMR2PE7Hbdpbr+njuA7
MHUSH4G8lP6DfdbrzPQxEMbABLWF+FJIepkC/EnX9J6loxifF2mWmPjHVjsDt1LLanCoZIWvrYxS
JVFHteDvQxK9exhJOyRe3HPBEHR8OwzwHsCukivkKA9Jd8o/Qa5IgCELVhoS7thCXkuJtOdxmt1f
4T7jSamwlJPfThq7S4/c+3GBsppgS5Qoa6QzjzO8a4Oud/aq7f4+PbleFpK5Ii9daQ6Ef0ykpPN6
OY9lWUm/pF7uPirZL02CPAjEv5/roAFiNiAXoF/SWPHvhgRrZrQ4qKxuWBbj4EOsgg6dYrMIDSte
pilxKOMQX2ieHrRWlCrQ6C+6Kp2Dyf/5n4GcRGemfUY6tLAfxVcXTqFC11ibI46W7XDlWU5+cj0y
8fV8YMYBku1OL6cUlCAKeiFPsAO1A8GCVNkNCA5iPwYW9b3oJk6VsYcKUnRGzZT1sYrSX3aUwT2T
nILaCQeKDAg/rLPGYcVJou//rQR6iq7WyWFot0AF76ojb3nt2pSJOo6EQp0ZZYnTG4SZmAOZbmX7
yoG6eAYApEfT4W/lRLhmgfiGGoCN+1iBVkicZvSV8ri4u0bd7X0lRQ0u5YUjgLiShYmHEm1/qn9k
uxy6+6X7iaBIv/+8HNw1ZuBoEiS7lg8F+0D4KOuK9wfxPVcp0qg2jSuhVT0CJmGBK9upDdRoKTvD
FmiB8y2stfWwWG9owu2Df6aH3BOYBRjBvPINykNcOGlYJmB94U6DFkwVcbPOv5qdP2a23O/PRxrM
u93CaxvKjZ6Cd9r18ZyG3cRtYTUnFAKf4I7CGj0AeWp7dRsBX35rd9vExoylv2snuu+Jeee/59et
3gN1R/BdwZMJJt1noypqkHtLaAEPhVwrnI15hhs8yp1KgyABLF2dR5QJxYt8IUNRLbTKQs1Af4yg
aI9kQO0D92jCo3whvt52e+FtEtojPHxMOYjUDyjLZH7QFhNpjlb7pggNHCWMDrFDLQ+2SFjRzZPG
NHjkfXq/wJCUsxCDIPLWa/HC3YEMqz5pbW/JlQSB0zzaR6AX+ibpggqXv4rNp7bWTIBIVGC0XfW/
6h/88f/WoXNLA/f9V26PScZGN589VPqNuSHyjxtLhUL+Z0eXDO7eMSStuM05B0cIOHnUecWWyHGV
8G9vAtQ7xCFZfLb77azUvrwVW5IX5nEOX0jk3sOaXKv/jjUIaQtTuq25GAT0GYlNMnmxqOy9qY00
IA6kmATVYvE4mY/fZaeWXa9ioXHlv1TQ3dxbyCMJl811jTfe/ioLcQc8SI5v5nJVHZPlxtvUkiWD
+xyUXsT32vfuweczBqEGaMAQf43Mi4T91qGN17nON8eX9AItoi5h2XFcObhx10kswVUKmonvqn6C
uavivPMun9R3330j9xV45sYjxgwgWNuI52QP/xccBnQekLor8NACBYGjuRUIGRmFQZSCOZFYlBEY
99bDCAF1L6bQQKkVGUvCSSa880ryIRis8c7XFyAoGw6p32a0yLFCnGRGTXFtPcYT7oOliuVt8JU+
7SVjYyDSCABA7/w8t5qYioNZINc519cWvBZJ95YiQjTngNJn5SSeM69GQKsmbyId3lbk9HG2g5pw
VJVr/D5GzPOFPmOVTivU5dtaviaXWDx2QOTDjWDVTIXSGslGB6lJDX2+a/zOyBgMVxq7lRG3rf55
vFBLlaTxCMO5zWVRsBCWRHyq2T/M0EGG6a+OZNzAua5tnT/bUa+caoReyFUN5i3y8F6yrYpxOErN
DffS4hZqGNYGHTD12P3lgs5v/+bIX2xkl7DyHD88jY0ydHfTm44V68rZof8+p+2sP0W4QsDZs2o5
HbLdygZzTmWMdWonlsHizfu7J1ykBpHDBiE5swGkrHdw+k9dkwxEHz4Efs43xlOmy7oQO/Tvpzd+
s/sE2d+3/nWwQBmK85txVPt1Mtxj1Z7JvM5KS0bUMZtw7mwqRy7GyL85fZlvXz1XUpoQRZpCV6Oo
RTPW41aTFu86W5YbeWrvf2t7lA5vvRrwedGwvZsv1Pz6n0vHx57jgPtlcE2erddGkTzOvoDTHuOX
t4TilgQzLA9hpEQOaFsc0RJYO9sWYCWMW3UUYVHPsmyadNbU6bWk/asfM9PnGbFMV42LsnbbjUz8
3HGdIEx0avVYkCVvQiXOXvKzBTfD5gL3z0O1ddOkVXc4aBuYWGljz6Tibhic8LMNeZEwzwqgkghh
14wAnP+JfOyKMCF8zuP8XgCx0W6QouFvF8OuRrkGlZUkFANJg2gy5RmhM2AFd+YNfnP7+1iy5EWf
gp2CWmzPfCQPDCdxNMN1jEeQiQ0hwQKFBAHoIa81EIIKdswVUfilM71xVWzVNh6b/bvVT8XFJ2mH
jB/n/w4OZCyTh8GBPlaDrbXeRibRGdnjf1Gi/a9+UVQ7QN5S3KWaJOLjLr9T5f53bGdhAvOZRiM3
zCCtkilaSHDVZtsnx5QrqpZviTK99DdqGG+s3MKlMdt2UlXG5rXfRP3UFWl9Ki8ONOhJTKg+nWWP
97xH84pdsVv1YOEcRXBfimP0Ci1Zvo5KV+TpprlCuOamzX86qeAuT+z9sTWvIN5pihZudNVihsDY
Q8Uewp6++2dpzSmpjyls6KC5cDSwhf8CLSx093gIAZQmEGPrWCWae1QH2T9zGagcERa+JIKLDpC9
Zl1fLwqTTDOcf4W+dJaOmZE0g5NVlXsOG6vvTkXDmpGdaGpaFvbzG1ESGCD6u6dL1yQ/QZfypYFf
PpO0oRKM/BR0TskHtMqG/ySXuoZJNncGUjhufd6D6Q/Tbl1VSc0RUiFyGFjebKEBJpCUhFPdP5u3
FmVqkP17mhEMYUzzZ0KJf5xOijttUvq81+90z74MAvqu1ubTp08axFiFDpoe2bIVOWs2ASw6+xqX
y8OiR5cKwmPXMjjFMgQBVcdDYYvNXqC6t0i/XmAURFvmqiKMpkHAPEgcqeoGftQ1NksUhKqkmvLM
xdY8/3t4KrQLMxHDj3f7NYk4QF5FwIiINvBqF8zOYa3QNkAmTkzMGyJcPVrddS9alNnpEmbmDKDU
2Vuo+RNN3zsy7ONDJxfG3okyg14roTlYfzNuH3s2MNj+3MI3ntaQ3VWjkK2mQYanyfCXf9GHQc1O
zL5PwNqUsncrv1QPbSQ1+GJ/cL5CekCsHKdMXIydXfx4ml9b0w/batrlNZ98Zwyvc7pgaMQhysGl
hvwnY/WiM3N4NPvTxPgjLiFi0XyS+uVXDaXTbcDZLs+czB47seM8HXg4T1DPVYTRO1d8mT4FNkC5
JT7Yz7OeWzPtqlX8U/W+/+lJ2WIxV/FcM42FiDVGqn7q3fld/+J6Ih2Wzv7Hey8/5T4Dq9wErZG0
VhTqLKMGDG2gwLsyUbngm0EAbbOYObj4RiUWsqsNX63LQKw0jgxXiX+cZ1JIHYg9M14uIS24HX/K
zRDfhYsQJzCNGwgySGO6vfGlFeSzDfGFFCmhUPHAuT617NUydiSTp8iMrooYpwuLJcylt3/OWNGp
8Ix/FBxwgSPJ1TG0EFoiPa9r4UNZ6nsCqXjG49C41ImT9+DYuBDFVXCZdLG2XJFebHKm/5xuJAQl
QRoVISIFtzUNH555KTZTIurXpq9W4ddDS46itPlp13LkajSsi752cBwLLvoLTx+Ilk1jNgw5LYHJ
TOg/gflgyKBw0OOcsuyB+BFCpd+5wO53GJhnySFpJ94gWr+W4bV6bcUALbXklTdgWq+l5MXhRCgq
LUrDdsS4WJUw7weQHFwfPv3+uO2Oc3D1C0LHhK3th5jaOGCsXluWBM1Eh6zwDXwTCNnmYf8tu57v
1NWK+6eyEmpHT+JmRFSw6OBzT9XxHTkH9WcoxKe54edQmy3Ux3jR17dz+Bj59IvWK2tvKdzaFM2Q
RS4ZheoLepZcSyBYeNRbcY7axPGX4DgtquCCtsFI3Kl+p2PRBBwirpNPzr5I5F41+/uq1CqLAjVk
HvURDnOeSF6kfz5HzZ/4b7mCPca792+Pga5Br5iUioRRbsfpe/Bol9vKA0wRD6kAJxboWYs6K7Ti
l/yT5MD/5ZHiswYuXSM0p874CR+V45i8R3+TOnYQPVG9rdYHOUVa3rQ9LcpJO5eeTwO4H55XbLn6
a7WNMr4+HFy6mi49hFl/MUiS8ySkrn96qi8wpAwNWOaPeCEn66seyHDmwF8x6L8pl8szFS2hxrJ9
pA/A8zkwcQMEyiT4WfsYLijG7RrK1UbEWf5xv7MvCsYes1oYbsXgACQMNh8b3SWtdfBfvlPg0BTx
0aPaucxEDqDUU34EumXN2z//G2ysjONmkhIGqbgjbuIiYYDPee7lcvJJz/0pTFv+3CPArNMhFFBm
1z/LpB2S4UMV+J0gZwvJEps0Iu9UJ3yKXqg+4H2unGtbx0H/e19PDZVeRfBDp2daGm5DwEg8sGJi
OsxPDrdE3C1r+QCcrNEh4T5MUUfivBad0P+vgujA62vQ7/DFikZaOb1p9cKz9s3hMUKRvccUE1ly
pkEOFp9pHuCfWdiI0HMpnXrAkO6n7KfkGZkf3erfVsREkCb8wEa2AZZIAkOwQ+3SbCiUGnxLcqi/
fXgU9mCTBQuQVwdpigmOm3LNFzvmHghu22t5i1AGiDDKkrATYu7Hn6Q8mXDDw61ukLL+33/Mq7Gh
/kJs9lJhtJ/h2aNjqfLDsZhVcOt3l9PryJXOZSqmg7k1L369QzWl2WW9l8dVMYGjSDszhgsdh346
ZqG0MhJAEqMa2JqXWZGy7jpaQ1Agy9Y5R064YirinIgJm0QD0fhD4AyJqTMqY3LX81Axzx43F/Xh
IVVWjuoQ82WVz30z4FPWMsw1aewjQFMkbtNXwnAydkSAkWkZu9emdQTaxSNcv+/b3HyEAdP42dq7
UQmpYiCprmbnw4DDtRIc/zHHhO+DERTHmYrgvNpuRGZEydHGbJDHIRQ+Ui82Flm6hQv6rv0PKPBp
scjzj2L6v+hYng/3c3Td0maEiY8tcln1FxnZX9qKmZ2n9P8jMxC+3OcXG9RrQoXJCsknNcBEGjg2
pE9SLkj8ULIA1pI0uhZTihx/i83hbGLL0An8W8IAN7qpkDEwlzl4alNt/ZFC+qFzM1XZexOnY3G4
Sl7iDjJUhZudlKycXH1cU4ug9bIiM0vJkMsRO5r9VVQrXq2UhgKB8ejosiQeNJsCi7jJUEy1HPNb
R97J5tbU/CNCzBeVpic+dhNMqf0v48anXtH/zow2JF1S8Q1KWXORPViVh/fH91+2ZUVvISd71crG
gb+f56+laYYHCunkeettIEucdAd41BdF/uUVQX7dfjWXK+h8vwLFRhZExLE37huc5L53Cj/yVd84
QX1g2Wl5UQmd03+rpO8Ti03h2rL/3IHDmbzamQUc22obW7lqTkT43RT5/aqpDlMgaBRyLCpRtGWm
qiZdFRP6LMOuCDWlu2Nlsi7b92qhAiKJ8d/cNmPQg2e2uSwBhrmB25mbGsw7nGvrpuu02OqRgsMz
Vf/izXVKXCS0fWDFkqeSBaMTo/60KdNDAruIiyQVlcMHgDk0gpOsCm4DNWE/OnLH03D4zghLQwkg
jDnG+/QKNya/r9jbXIPChC08HbAD9ef86XvgbwxdZ0Th8akWThyIaB7Rd5BNz8jC9sgm9TY9cBQ/
H4E1yjJhT6cYldZOhQ14l3LP/ZAmz3u9CMABmdnkhnGaBPjLsoEt2TYxr0pOWpnUlOJEN/6VfeQf
G+f7yJ0gpacH1JHTUS7FCz5e3dIqCsO3S76bGMyU1OulS0d/essVHoqswkcKvPP2iaFVNqwLgEhj
eiW02+yCGdv24laG1Q+c2ch/NQ0J4I1JUvaFuXYAuAUwskMnT+km7RULhGzxIilYVRgFLkrHG0AM
OG3QKIL7dYdVbYRTXrV3EDXfjlu9ZG8gf1GqMCNji923eXT6bq1YaoHHXxjR1lfL9xFEfbHEVC3o
aGLpt9kbzypl6geE6MOCunmD1aU29gMvc3AaN0Q8YojCdcoL0QfsR4ZJojfm0CVYufrR0VxyGWK/
VLQdsugLWr37jTbu58QqoYkwx3SHxCxk/S6j2Sro6bX5sGsdUybZ5wrCpABqdOE7eoB0VuKtsi/y
EB1LpuUUXn+TjzLO+Hev6L3bhbhcQtgubYWguzA8t/zaGMqA4HNUPw7jWO35WI6JZ3RVXpsVS4lb
rENC3eoIxLTzCA3BYPB94puvzwlFqMbjQVQxcwaJqRGH1XtY57xAt4Ukv5n2VWPKDitqR86ejm9w
9gGiKq8QscyUWGjqhT2WLHzQCEyAKUwWN1v7AMqsY+qzX7G5Zji0tFGLvE0p5/FFYVhJpV9J2uak
HTwq8l03+vmmZvCXgVvR0U0qm+Gk34S3oAq6n0jhMyrt6E64sqAopJEvovwfh22PP23eZzMalQC5
xHsxQEu/x1xNTdVvJ3NtmPG037hxlR1ms91zFhEVxgkZiEAmDuujNPtrddBhrz5PHDqppcjtOh6C
aN9t9HVfZtaLBLd3GTIc7BxPTliMO/ECPv6d5B9iazbYdl78BpJMsVx5qTUnjHboT+x6aXhHuV68
iZiFFsSyGN5LC0NnKUf1SB8ZxvpHZiKsUmpIV4EAzQqNCRjzPOeFTvZy8dhdJGjyT31M2glqcKtc
yIK8N0QKCnWdLbbkWseJTwTOxXIhK9x5kx8+Kwo9t3mGncJCdeX5XRT/Xu5zx3c+pH5gemBzuIIG
CuzceGmScUXudOhiZV8TrMLet1oOUxACA16/xdOiiHFKmtUxU6nKJGJ+flUtBDBm7j41muSIgIHD
cSbfamN0VFZvFNaWGZuMkRHMOjsNTcE9R91KZzR2bqttCc0ohIMMUPnyHA1iQth1Zc0y9ybnDvRX
e7eDnl0mEzWmx+RQ+lS0v4Oozt7J3d8/HZyS1d0w4ZoWtx1li+5se8xhAM23T+p4FAQLBCzNZpHZ
//+ywg+cLuwaGdYmB2zQoMyJzzgmTm52gksWeBR8VEHXgJxAhRi1ehyG5nned4MIAgj9dXnL+fUA
HoomyGBEwngS4CUpHlfKdMs3NQGerEEaDp1IvxH1+gl1EHBaADrZmmWJscTFFak7nxqZke1inQog
TruVh04SZM8IbjnXHwP2TATViyAC2XohCVA+5paPq4W0ZOqDBU4wWmb4WON6TXx8x1wMxVEm12L3
WDKZMAEBgU7xjS9kmrCD5ogV56kysxl0UChqljg+zX0eTQDmxWvYvoA8qPgUdeYSOH4MKZGzePab
3tI4yDTu8GRWU+k3L06zFPkZZaoTrPBazqXBLphWGzx2VSfjPZwryGWDdVro/AMFYF08x1wFda01
TAN59WRB00l8sT0HCsf0mVdNEYe7kl22yUwFfJxBj9QmIxbaFLhIHL4Vf3baD8MG0+tHn2ms+wsb
mYwI7W5MULZCfWNFXu932hxps4PwOSqnhGwWl+QBSyIxcSwohZsNuytepQWCepK+4msSWTI82Y4H
QV9108HC/5CfrYtKz6X1aYcqAgwuh2noN45OefKK7whIK8qvq5exH8f5rBdi1t2gMRR0UMIwK9hR
zvtueO3w7yx4qJv5rPRzJNKmMNxfixirKZNSjquK3kZY6XrstxB9fswJJtUqGvVk8BWr4H9K+NB6
VtIUrq9CuEzY+z7Eo0hNhN75cKWoZDkbbJZtGiZ1qJTZjPS8bpQOfUQe3rh5yej59NEfBRMhvpyf
cI87yM91PpAnJja9mgzhCanJv48fUl5a6FtXRvzjMYd1NUjVgppuZScQ4xFX2Vlno0SYNEYQuMbc
8WcfT934iWVtLXfyJhbUTPNfiinCUpd7LCYDyQco2ZWAVTLK042hYbonfv9XuJ7XZBE4GEFR2fX1
/Q/pnc0l04HQKgRdQFW0aEIpquF2Sb1BHuwm2+P18ctNdLfu81Uf1ToU74HjqRIT0IyC5Zy8R7OS
B/zJFWcBLfoBWdUNC/Gc6tGTSyGrfkgmQzKrZimXS+srYI06L8cRtFghem9REwJSux1R+PLUWy84
tpSgKgGjlgf6I0wFE8SknyfoC1dF1piVN7Xh/+l6wo/RW7ukX6GdXEb4xFWY3TaEtW08tXFcJKPN
jut3KPBRQyP1e4NJw2sY/q42nzz/yc+sHVfz3qHNs5Le6CHOheIVVcLWFrmyX8SUgzizqY49B0BF
sYXliFAOpXHaOyAA+kxHZCYT/eBTeAhg3HzEi4WX9nAXWU3F6MQ121Hl3BD8pm+0CKpHQXkvTIVf
fIZo+X/7VCh4WUh/0AUh5GtemoOlyMBybcG9YpA+p8iughQ4YExZYmrcT43+Ujv1ipREagr9UcgI
nDfHGt7W9jDb121Fd6fUTsiRRaJyP/O5VmSghiNruTo4MXH0LooXxcHTOJ+nJmA8K8EaGuJ49Tkq
0FcmYUMDgew45OKZLDi0gHDMeSy3u2aDKxMj6deBoVgUaw97OUl24WahF60T4SCXxdxc0iIqZh0T
pcMVvVv/iQvYr+gh19B60WE2QqnHWx01K3h5w+Xb74rttSRXbOmgWkz02WyFkWXi8jGyuJiZkd6c
tIUMgksru/o+pxizHzcNG6j2b0CBMLqfMB7h2yNx2ThHHtCrMU9VnCEOaJYgtGwh4YkeXQ1mLV5c
vLqDrwgxZo9DOxW/e7s0gI+WCitVeQmPabYyPLjJthKoj2wn9yzpJ5dlNoboadSYaxT8wr1ePZ3r
11xmnvGE//ij5Oeq2Y297Kf6DOafLTUBB1AX1eNhQqk0o8FQ+uOjea9DRvim9ARufFq3nFW0OCly
ipJDIerj+HOUozq0S2kZXPrHZKGjxg0wcuwbbs1hHST3JWVZrXTNXCA6iIgCku3aRqgmNuBLJ6IC
i0Pd7fozxBQ8ZBwYY8jjkm/b2y60y+2EGjFhhcOWb3YxnsEVF4eO36J075UidSKVz8wJeN8qeROO
ObAfjqnpznLjLgDiR190fvUevg3AHGy09saVhJuhYRCL/fqsD3jY0dd8w+RVV+EPwjdUNDo2MCCY
V5WajwG6WMwEz/TTp90bxN8t9EHTXFOHmQHrLzEFvmDLeW9LpyrebkLQeLzj71oPb/FvxuLt/LNo
/z8IliodG4nMa6tNhmlsBJOGw0Ne9/iyrUc18/mp9PPviNXCHaDWzg5m30ZocYImYBQyxGj2DcU3
/TLwX7b8V2yDeOQ3fqbgo0FN49WR3FLmlGCJsJMzezVQ0FN6trAq9xXjCOhALW0LkMc5tPhVYXVP
gALPi8egcxPQUy1LJD63cvW53JEh5bdAbm61OdxLWXeKiJjq9sSFCrD1uqxzNj51dhQ+WBKerWCj
Euh9CU1ONORvE4HiwekuFWZDLR+920O6oH0eGvmESg1z546i+uw4mbnoUAP1PBH/PRkmyZnafScA
OXmm/Wmg+mZgJTJiXoDi3fgB8YVa7SEB3cC4q5DXcEqyNCNK37BTmYJVvHDX3zhQCBa2PY4Apikr
hzxrvN/WCE8w6CFmIdBLcUxUYuKZ9S6D34Bsd9wZHEWIhRF+yz+2ChENLuQu1ZCgto5ZcoxNvT7R
WIkfhV2I3woNZvEypbgcJC0E5yImeuDU7PZ51a6RfoVb3b+CkIKo4ziwjndQI56JhIYKierg0efF
xMCv08n3/CsCpuAiFLAPdwCvSgm5/7hvgLlsghlIbAyH3H0EEpc4/rcus56uzMEml8vez43QyFTr
km3AfyM66MDp4q6nl+bOTZcsHXXhtDG9i2kH/QnGaInFcDrKXwLyD7cF63fwrHZSAx9WPK9Qe5bl
j7ylguis542wnekXZ+Qbh+UbmijM24sl2itONq2jzmHqhxfwUNeYKJZtry/NDhYw+2c/3TCSS4NX
VLtdtvT7pk++mqjLoMq7qom7u/CurHtnfYUevHWSEubyA3RfDuONsMUkKtPsh3saGpX9z5iP9XwS
4Ug4bFSby3+SR4tUy3O28Q68ZOdFdaAK/jBkrtoPDh8QFXiiUPkQT2O2aK4wnp51pvHGncmFXPnU
B1rgb0bMwRa4d++c9DXZEfDfP8PVJRLeSbSakYo3VtJ0PjM9y6eluqup2ZcAxFuKpR4569rRrYqw
MX/LoHGDzGc0t3hiDaVBj6zdUAyL9JUWlEtrSH1uOOaY8c/ZrbCdrg2b+JNkvk9ReeUwVc62qw+L
MiLUasP8ngUx3TGj/20dMkJXgcdbOwGHrXngEIwzKxl08epcMGWptbVuRPqL9LLhUiddJmjjKxOp
kP2eRG9s8tmrqQR5jo4zXcWVKkGpf0TaKwFTtRXvWspXStrgHqVEoVPlTZgq9LNk+eWkmloJDW+9
3/oPR3QChkcUdgK3gheSwUqKmz7gvA4QF0Gjy0VHq+fMt/nwMgxhOodFrrA0LW379sWVOUEEoJrw
XRC1IImv4Djvb23ZgwekPxgcy4GEQ2PLcCBr4Ch5rlNo3GTkV1Dd1zh/u+2TDwNw19GhBIYPfvl4
QhTngghrED4opb2gllj0azHa7luXf6aH6XEK7rsPr4X2rmeyg86rVGErAdc/6UdG2uT5In2A6te3
6JCnrteWbj2LsLqgMdU5ymjDczsVtEF7lFXCeiKOxeAwqZx/Kdqj2k+qQ67XM2yFumdrAsslUq5L
WYvAUeKSQMnAFaEBBBK7K7QWNgTsZW2LN50n7ZSb+hIBtTZrZBzzL+MO4Ax3Lg/XYiW6vVs/2IzG
ugMy56qNJjh6/vZiSmvIeRUT2Y5ZZIFmdFRixc5i/uRgYTN0Z2cFW+ppEu9ygFQgHcDQzpoJtQrh
WoXDX7aPQfZQYsbySNuTu+r6qNra4CeHja2LEWeDmIaDkWUFt/Y45XMBLY81yC30Acn8bu/M8u9I
ASPDgXcKfWknt+AXsIakiH34YWy9+N4NZ8C2cFryS7TohcDRjyjciJidbpQNc5kZ3IQf3n9Ug2pl
dmKXfRIZxTXqXMOyOa5mkAHPHV19BvXyNhGZ0Qz/EqU6ZoDt2NT925xcI3lHbDHh+ZOSKBoNKn94
8FSuGG/QQwBUrpwM+64EWBVBYTqWXxwnNdxzVxfUHM16LnRgjdXdf8cwFH5UrZ0wBi6KF1KklvjX
HoJxq/fTw8WCa8iMaNeIQ9ZSF7OgOURuX0CZOl/ktJr0I9+8mU8YbRKFiu1Lh3j1BqBlYUXFxh7J
dzceQbMi9RJ7FTl0p+JzI4H9GIhmGClLS2Jg6fymIJZtD8rFOhzLtcNeh2SgJ62ZdHPk/Dhv3ybO
hjIN6k3Cdr95YryQ9WmoF4QPdAS1GSjeP8ZrD+juCdXzj/BudIuUzC2oqWamI8qLSPISGbcRVFkq
wTXIFh0P4nQ0389N+6D/S4sk2grqm6FPpFJ9BMqgFJxrxtAsKkl6wNv0Ssn6G5uVzM4G3zciOueM
j3XmUzsLSXLVQej23ehEEE4sHYQVUM7AMVquNJmGDSxpHZ+9PYJWPaHIYsrBXb0WjgciEFKIG7/1
ox1/NCjobX2evmbAyW8nTq3ndNkqE7D2rGBJJ5CW5u6m3Gpyf3cmIMTLx42Jh3E7VYqT5moda5NQ
hpYovxnNj6qbBVP4hdhZ6KpK4SpiHLaNFZzALqjLY3xEkJLBe77C1yore/bHn3cX7MZMGkt1WsfA
oqsC1sPRDEiLVJ6ZyGdi4LOkcXr+yWVAIB7zeTYPd3y4/9os682TsFWptGUUjXU3+57xc/5DPjvO
IH1JosenFuZ/nrMOU7t04TEonQG3tJKefRkKAeof97a6QDD/bpDZYVV6iHAf5ORp3IxJIBip0bc5
pBi/nivMKnuqQeoyCCYwFzUp7Repm5//9UExK+2oPwugknTBwQQQdwVKKHA99Bkt/iz6f9FXKCrx
t5BuRx1MIM6m0Rtwdpfof21inzoUkQvurMyHiGXfuH9wdWJq4NIYej0CGlhz1oBziv4ZdfuaEMq4
CH2CchzH6RELjFnJrJnnDyG8ABqHdWJsq5QJX0i38rrBRn+UQKlMtd1bgEeoQ+QLqfoHN4RQFP7r
D6Qq+Ssueb/ASTDQWFIJ/F/XRuPt9LMLMPBy9vDKUtaVEjKVrce8kVsNN3PGPiadKXN9FZA1CVSz
CmCanHnGZ1OB0aswQzuqoEeEwSKItnq6Vx86aFQFyKP8oDv/05ZdckMgJfUh2VEsZOFBWiXcttar
MGtbi7IFT0/tjDVkNey6GKpXlI7zH5Ol6m0QD4qMuRSyxXT8eg7N874JrQZUsaQ8Vyv91tbVhniD
U6NudkA0mTE4rFxJZA11F2arB3yRNQbGlFAjs+k9JA/Y8Pk4LC5lgaFpzjdDfqxJY5LneBNram5l
lSzVvPBpyWstsXwCrPPj8q6rpDVW/Qd1raPs1m2oIBEks/i06/v6FSMmcnUm9vqgjIvNLm9h12Q8
5j9bDcTXDcgPplV205Sk8jN+hOpw+u3zKJ5S48ur+Z2dhzfInGdwkk6NgAn1Mz9gtba1Jj2qVZrj
F6JPnxenxvCmvG9QOpqtLOuyN1rd7Y6XURm0gYutWQAKzhOrgwoElTXfo0yf6BU0sP2LSM0OiYiC
8FteMyns2JB/0TKBpf0LYbIc1l2nhJbpseTfeKL4LWirDFxSKi2h+Zpf3JdDwOAKCBs7GQhyg7n8
BjgjLG5xsi9rhvJIvytxUoOuPEpKoSuFU0f+XnOyg0KXzpw8HBTv0xF7iZtzuTOiWKbFukK0XgcH
V0A+Q5q1rPpmmdasA18g6k69Dyh900Z1wowiKzFPg+U91jbKE1C7MQSzrcVy8MvmnDvwrKEA7+Cf
ZtVBXcQQi0nJ7vCaDdBttTFJTVvT1BVd0reYDfO14cRBudvcnBe5xfiHcJxOwX1t+B4gTlT4hCqk
smuuBPOrUtaYADjOoFvpOByMqyu+PWbcUwac8sjG56q4XCMngGr3IWU6sRx1a/T3dxCQFXkKdBJq
pd5doNPEmCaWzMBXB49ODzwjA6hKKBBgVEPacWPsDdDZGAKwYu/UbMixtvNiBC0RKvgydgrGkQtM
ieq/lbG/4UYGGrPeiJSvt/pW9Cuo9SvFjnu6B/ugtSNM9K1dlJvRUG9vGCaxoDJB1FGeTVu9RFKk
lSkwdBGVf3g7NjGuS0BRbVirOCchIXGTr8IAFfo7mZyPVfhnuGIip8NeHfVCMlpPQJ5gWz5nuxG4
wyG/EBeB0yJujXz0siN07sTp6zRbZSnG567dIWqv3zhEASPHn4HlPzXivwPi6O30SUSNFpEW6aXk
oF3SSUBio1yNsaItuP1j/C1EPqVDcQyLOufS3LKSoplZebGZ/6s6aI5UHxNRAx1UbyCI87WyNpli
1Ixyot5Qq1qTDFuxVB/t0X1CE9PEgEhtkyMVTsFu6fEO+cMjOAtVkj6BQQ5qXSGDxFPbU0MeChQN
p9Q5WGFpJGLiaFvLzubDVPCG2aw1fdW3a32xIAxVvszZN0ShILUxMq/WzIQr6FDXkD1IJ6a7Ea1N
r3D59KU7NmCFTD9BuFwKmRMwZMWfeNIQlIM0rjP6xldtRXkYMkZfjEYmwldq5AH5CLGMQO+OLE/R
PKPQF20I67Mui7UiOy2D4yKEP7jxkZm50QS+7YLcB8r46mYa/8UnhEaCtZcRLYfWnWVMRXZRUUN7
DDhKp/JBZnAw0f0qFufrC7drrOFBIdMCEwY3iDBA7ZeZG+5Ai4xfI64eO40bLtqiRDPWNY+GAujY
trKErch5BvzhP7AUigkKdPUW+Ht1mdqHERONDgb7uXjm8UadKfhDdOeoGaQ6mrGCRfUYNqhcLOp6
WWefYG1hsVx6qxsfjk6gyYqB0rA1S5R4iau84UDQZLUb+QdPG//HhbqElegm1cVYMubyuXpaW9sB
k4ntn79GzKDK+mqAspN7uFfORYNEqGAEVEKje0zjIiFAX0IZo4ifM4PxjxReE7mN5xT0NCnu8pNt
cNdbNE06UWeUH/ag20LMFkeowdwR1HuEYJiwEDeSea7xocJRZES01Wds27mh8cS49oNFdSyioNl4
w1XIS1x4iEBREBI6ghUjpIzOje5KFeiwUMSSCpczJbJewDW4KfoROcsNK80MgSfn7D6DLeFeqnUU
zqObru+a4kJtJMUtlT7EogSeHLaqTvE6WVehhRaPOpSGmOLVTLM9W/2V3aLpdl97W+4T3DzcpkQ5
tEFKZeHnrzxXJSK8eSMhC+70G6KVKpxoWUSNRNBNw2ZST2+p9GFtylI2fWbyqXIcNPbWTdbYO0JD
pfeQIkAppuBZjH1KmpfEEL/wTpXbRGbMq+t0rGILjo4yg+d5//2T6ndI0gtvmTBBttm2JoBJXJ35
BFKeZPRoN0g2U3Ukh6av1EkGsocnW21yTLZadZsTpGWnc4SEtjKaYKTIjb/YcMCsH40eTWCnbQSK
m20yhWZsiTsE7lgbv6ZQuFbhvarN+TosNr3qRW6viPY7hUfl/czB3Cg6DnVpv/0jBz07kX/BCLjL
AW2OM/Yv2PqsbLCQJjsvzJAmSHAfpHFgClAJEWIhQ37puwW0lnk2xvuCpyl7myc969VSrtCY2rBo
zESorTOP+1XcLEy20rSA8XKrQ9BQWcZSDz96fNiIlCAGkVWC9Mp+pZTk8I7d4FfIEIHqbnILGzVs
DhVX4ZPrT375cr9VvJMQF7qQTAsTiygYGMT/90bcQiw0wSCnRxGvKf81ekd96zNGG8JWkNnsh0Na
/y8M3t/+uxzFnvpWfn5GeiI4hc4ySfPCzpOX/ZCvRyIT21b4fI67rha3xPb5yfLOIQrk1LmHpzyD
eYUk9QiTjQuqiNB4EM4cupSBEvrecvkTK0bRnWr4YI00lAMjiDGF/SctNlaCjU+sJSwPUbOM2Ipd
ovVn6Y2DQXxPBzE/Gdl44oN5mwjuUdQxcptQX4GCAJe7G4RlpYl5ZtRqWe1akSS6LsuZTvueA5EK
TtQPYsg0GkQTndAVStqfoW9BktPs0c6aAxKAgGgL3mQfNJu12uBhaItxD727JBrgUut+6zNIDfYz
g62/1o0RfsqOcrVsHl0hGdyH7W5u2q0DOD7P9um1KzdbMBdbZGBcaP/WjS/ud19e8tWvukjWb1X+
f2CFdcjoT48lW4MxZYAhUV62as/PU2FJH8srHx6ZAMIzOvUG08qrPxc9lE8P6H908IKBjubmHeFM
2OSzNWpnPktAMjlqPstWdYObHoud7sL5FTmusK2TrmFB4OKdYIXvd/Bvfds9rWDF6QwxzBSsf4i/
Ol++oHZIbQia3iVHMvu1Ci7+7D8GgS1cAqWXk5NaQ2HlyHXJsH/Ht1qcUoVjJdBdZrHbE6mvJ3sF
/UlqYPPgzkgSE9zHzTMx2hnQ0ib5JkOahwigHuBCe+UCD5oGGO/MG9gPezVgoieAaWaoTY2DmoCR
MS6u0xtUMY5U4sr2qwT1ZslUTExLH2gtzudiDL6MElexg5geP0KMP7eONEnIqoCneg+yuQCP5DAo
iQRJjrO1FkHIUaKBG5+fiK6jd8pjzYQRyEKay51XCGBvxrKMpYzVzoE30UptdUP1uF7ZmoH7P7f8
SmwVegF8XbG9jE0pZdI+Z26/hoCB4sgSBhI3zJkPurT25V3eyUs9GUiO/k8jWc+qNbOReUDnMoBO
mbY9j3Jp/UThtHjwdOfHUuUydOY++K72XzJsfEhap+95AcG/PORYVtQ51NdLXlzU5kLVBR6Qgo/M
Bi2jVKULGf7VdpVNPRP8FcUpY8f+bB9DCgmHQILHA+JFmO8ZtaDF0wKyfTdqQuBHYhVOlDrlsP0v
dmHUC1hBY5dvVLl/fr7dm0hOTmrb+21x6at5w85MDbyLP822UewDy8MC+k+yFoZgKXVlpA0/hMpy
cBQpO15fjL8isIncSuz+17ryjRS3nXKwGBWqaAqGyiOogMDy0R+OMSqsIDOrre2eJsXxDhHmlzLf
UHMFk9pjk5WLtf96Taj6rlEqzyCWobbEtBApk4tWnNvK9Immwosqp5sckZQkpXHLQaRlq3SWscBz
/yVtlCyc/JMiIBM6iPBmvzwwZLxI01Ctt/M4HtXaqQ7mmK9Y2U8jMHdCKvor1U65LTt8AmD4Gai2
FwCRwUG1Tz7excd6TNLH5TOLYvIMVKWCGXGk+aTN1Pi6Rk2v9f8o/FNTcyT4NME4/59WWd/8kL+d
sTQFIOKwPRTNmzULWpjYX+rFN8RoRCvEFeEPkg4Jdezezpd7cgRVAFKBjS20UhFbvSJ/+drPJiEF
WB4Sfi5mb58LxgkFYTEdPeJfCxmT3u01cEhja0fqY7nKD0oiWO7Jh3L+rISDA9o65qlr2qpeAvOx
4bN9yufX0OHSOC01MIrIKJnF7L/vCKnymsUVpMAxYGZB/NWPlf2egakfBDyH/mm09lBaODqzYxFb
/O3NDku3pAES1ziy0ObgLf0zTpNqqBspO9XYV47eAjOuv96koRCSQUjtqMAU4sfbdHruXRc759gi
FIFPmV74ivWQ8Q/Bx6CPVQzyojyLm3Qw9beuCDA4S/3vj1484m9gaUjaUZJ9gkW/iD6QTQ5gAD+c
24bUdVPbb0Dbrzzqz94piu7hxByMYjVCB9AxkWo5YNYpcP95xdwaP5cq1U8f7+V+s3USZ5u2iU7C
UWI+WNWgGiMQVx5K3/hBtZtsIDEMErVP40X6KY910Jjh8HB+rmpRsJfOik6SRxT99mRFhGZ1/Oad
cxim0+lSt9lIg0K0l9awbx/DBuOx+Yit5DlZ2tz4NIjXuAlN24b2quMuRplUDTZjCeYBqNfUjw4u
1ZSjfYOKrPGsIOwNKXG/ZS1VIQEPcXxSDh7p9dI4mx54xsFSeas1Rya/ue701PXX/QpxsKUHKEMN
8H8qXx/dYKXk5QR8SLw5c1e23K0mmU1cb57U9Yt3bm3yndNyqE6H076AmwxbnBTdCF34HIe0ljfT
8Y+ZJdw0+feJR1tBQs7sJMwH1VBN2vz/lhtPhpC+vCaF1slqdu/3BF9iLvinsYntUATaPqcIrQR/
TE1KffR/dGIuJULzs4A5ULL6iwaNX/phxcgYOxJKkVGNzu6h1ofsO28Iu+cjY6vVyS7IAa3flsLC
xpm0xkjKY2BrMzRdVo5DrmcLXwiEj/iNuxeQZBz4uRd9Vr7fAICLCyhL1tSHoFeGGXMhGQeH4ZH4
LJVvqRDKxQCU0fNug77cUdHgb2ylkbGB0bXuuOkwsApsOgPdItUliN4sJxcV3S9VEtQFEvAxjETo
jjhEVItQrdUAW9T0j2AcAwfucGeToio8I/XhlvTI6V5cSNKOWXTIn15iORCwS3q0ADWQrkETiPcG
vQZN5N9O+2rkEbbaGeNd6T+R27yawVJOMlRUxl4USQcnFAEs3zDC69RJDt7OcQ1zVvKBIVIXyL/h
3amIvjBGXpb0atfMzShiH3YlMG7AeUqs3pQLp5QgsXD2Jl5pwGgRHnkguWMwSEUUWyOF0yV6EsJ/
UP5RGcoxH/tQJsR8n4AP/0HYd74Nc9SD8T1hCDwwLxGGLhLE8W9U+YB8loGsXYuxwTTXu4d3yYpp
OH8MW/5dIflTNX0bmEcbnUw/VDExPq2/Q8O08U8typAvCbEyVmaVqtU3D6/jSRRu7cpUBQd1blsO
Jsyt1P5/fMAaIN/cj57iVHWkDEQV1sIxqg7utKGZsJlyeuCPgst7uuCk6uxUWLkZuG8UtHoPCVaH
MrznIKO6EX8diOOYBQbDcyzpbUcq22q0e4m3htjGIlqUoIsZPWTK2kczEHS5IVL1jA3CMcI0ikKM
kwCy8P4kXu5tGPTlB5sw3nvxgkcvicMcDilIbPvOVxod/SEoo2nJCn2UoM9YoBdRa21eU5BYN8gq
wq/NT4o+OvYMWJEJwQx27dHOLc++tpC6Mf8weIl6nLv+QjhXa6QyWlxVjxAlpjuvXmCwABCsT0yy
ctXl0cmA6jCaPXLZ0IQgv6piT6Gua6yhBFwar1njOlZGFAp1Kvsr8b6SQj468V4MFKFBUylHsGoM
/prixhT+eAkpcbLFeM1xTEkd5uUpTR40lgPwml1RHQt+wt69VdZWqKVUi8+hgbZzCfIBNYQjoTyy
oDl4GqHEBnfjE+CjQyq50pnrJXRFcrw3SvX6Y4UFsBPIq62tyZ/E/+UgDs7qy6rYSxKLww8yP4lF
/pO2WeHFS06/+TQVidjvjotwh/zbHPYOHrKvyY5c/QujvaTptiOED/GZYnyBHC0SLhnVHfDbReTw
He8PAmtMxixlNIcLAtfxw5HjSzdjF5qR+jFuSRmW7tkZP8vxCqiVcpKOQS+2ZyOfge9LOvkeLniW
/SLveHK/B8gDTRAfEeOMP9ogc1l/BZj7RFGCTnpp3m0UXeSd9b1OaHvhkB5h9d7tRzmc2z3q7bKR
tGT2w8idN6coRMaAGJKbQWeqGos09DVp2aonU+83qECmSYzmmrw1s+GpJn6i//jyc4xQOZ7vTLxH
N8lAC5XGleGYS4muMb09T50r4PAsFhEFBLW13Uzs0rtz4C2HLL1gLGFgOENCQmoXMyFqAt8Tx5C2
OtGe2yb1eJZr4MJUYAyBYMTYeTqjKPilQWfc3Ti1+CeLmerpMOavBbL7Wt2pX0v8GUel13HhH/fM
OkBBjpjJ/GwdinAqTSSTlmIVxArw+eG1qLDwfUMPGIlotk+PunzkaoX65Tc6ipi2TJ46rXbUACEi
OzzTRzXZqsrnRT5VOES57XskOrjqiJYh3bBcbTl3vAYJNVY1c42BkcfsLNXPUHcwP50s7SeU3K7y
WrjwUMMPUlXc0fHcq+ENMa9iLNDeVFzvL0TPdN5n15LRKffRzQJXEvukQFrZgT+r0qGIyS1zh5H0
zwjomGznlqQccnaNO+a5JfCF4jZw/kvR0Zd6n7xszrNHz8efHvKWLXb19MUgj0yCGjbytVpTCHHi
/5OJJtSp95bAydaMKePsSTjCiD9D65XJKZvSeLkIOEiE11borRGXUOcdqxRLi7YE4CCdv73MK2Bv
i6yDlVdQEjAskqNm89n2ZQxxWsjzCm4Ym2sF0Ji/tN+nFzOKKv5dm9DtbH99Y57oMHW59zzh+K+7
DLaBb8M/ZdDyM5nOxxOY8BXziwI8ixNqBwWaVe3gMuF2q9w1Cr95yQ1sa4I2SGDumtNBj2OBmwR7
FDAYu+lgNapW6g0GcKTF318Q7tCzfTvQlbfRSd7vb1MWHMmqmn33Hjma0vV2oRmec+d4ZAqYbykS
jJPfjlwlY2GirMh/OtRjJfXsJvSlhgpVChqcnrC1T0ei2xsgfVry6bxrbaBXKa6TgCKRzKiIrSB6
k6XHIegEhOrcLqOvWFFvyiHx0PY/EMofJBhN1X48vPkjwvgT2bcFg5kDDCNgv+YLyLJQCX1vsT9B
Wq8on0brxJor5yhU11s48mRYrsvQ5fc3CA+QcPgPGI2d9BOmPOl8kuEvQNMy6QReTIBms98uyZez
7xhiUX/IFCEY+Go+aybtHoCufdlpwtyAhyiQccMJt9hUSUnzBAMUzlgt9SJhOSirpA24rwA6Ztnb
WsGLXa6Fr+nEO/H+lAZwV3lvxKIWShVi29T9t9yY0gNC01/5fdMgvnjjrsTg0b0FObQnWaC5vKp0
khcHj2ngS7PWsNYmVjZNMYeZO4O09WouEsIOfGYo558AKLmJ7X8VlPdKIaPuyBsTQPyQxdrJ636J
L/5AUKPS6XXBj5VceS8UePkt1KX2LPvMcPl/e27PSmvekT1JoRIoPy573GyqczhQzATg3nhPG7oW
wtoDyoNBjTROJpBSnZ+Z8ehX0FgeOsB4niRMgKMOP1CJBsirsft/LxHv1nQiEOJmI8PvNZu4xSAg
wfueby+1ZuNFz7cklHG5q1SA9GaL1DJR2c0dye4I1z625cOF9y9Rz3dxILXM+PXWJgy2kbO60nf2
H/PHOK59kvKRseHmSE+GDt9vzLChJ31leLdHarJ1lk60/oYqQAp7iC0y2tcA7wOX+H7HLcU9qUAM
t7pZgNtyr/OY8AI2+4u+aehknFpqDGb6sQV2KocpHFe8uOCdlc+djphPyeDB16FXQ/2CzrB/QDFS
WyTaKySAQG0vLLOp05xifUUQo9LwD+nmU/LraAcH+nK4Te6lcB+iQGazLFAc/EmlSn/Qvervv2Gz
af676RjeEiMrrtzDdhB64N+PhnxMjXT4rKBu8OxHMtN4updkLR5Mqp0xsYvnnWtwyimU9z4VDEON
eCYsa3y8m1+a1TogYr+cg4yH6xU6yrs0nvOTF+2Abgw6+w9R7/hh84uwId6FrUaEpTevoWHku3iT
6UNeyhs1uEK2a4pRaJG92VXCd93YAGKH7ZU0UR1wu1hDoq4nmqbgnENVYlnmO3AAxMa66U6uVQq+
cS4lf90x/atQAGH85sJ4xwzByaH/BMIo9Shb1C2Yme0LcTSq5WXK/OabqRJ5U01sHhChPjgpctuz
iFLJFc4CYykLLg9VjSo5jgBtafILvWsNiZbJhIExugQvO57gojYFsDWZ35L6/KrERTf/olIFtZEV
bIbjgkgvKbzYaXTk9jRxlp8rU75/cMp+Xj0ODRUE8rrhcn6x317cJt+9/4zADrPzX8aCCX0ECgDZ
X7ZE8RE94S7Tz//OsAnHkeXTiT4tZfqHIjteVE8q6X/tAU7AVs9BH5Klb836AtD2MEi8n0m7W2iI
ZRU4CbwlD9pS+jWWfRzM/XI/N+U39N5TbOfKL/+p6Ro9GVCQvSchAoN3rWRKxEaVonWFPnJzh7pl
4yIL+Or7+xIOGDQJDkfK7cOTCVS00lnGaL5pCKHBUU0yv59jJiRcaxpRgze+8yHg5jG8Z2OC6oJw
SQ+gB0TRkcmTBhXXo9U3epsLJvkSOcbGVdI8eDNGYpvy66AD9bYR/8pDlws5ZAx7fxvjwdPwUZ0B
O7hiJMf5a4bZcKiM6uOzhzTRdDQRVwG4lixzjvdfCMLUrLpWMtLa28PGP+hlkiRxLpHMTV6oNiV7
QqVsu54LQgHjz4gZWz/y0RB8ZZE9jgYXuiwa0NQKLb5ZrOFsF7QZMFkO9S01bYxA4A9u7WLxosrN
vLikBRyNSEFKjBeHBits+reRHXeDtWgj3pLvCDJJBUbBMa2tkW9zvbYrptNcoeYmJbAQSJIZLgWX
A0V2s3fwo8ebznwE8TZF95VD7qwVTOz3Co/IWQGCy/RG/FrC9/1ac1iIIYuzimzdkLeEBeXIP9Rm
gi/FWCnAr+69jJNWfBg7/Mmsk5Qzit/BlUslmswu6ttUU4Nxh6Y2GvgzIX52DCA9NtZbF6xof9Jd
8JBAbQe14VtqZjS7VvUCyWSqyxvf8lRGjE7mYa164CPBC9ybbWBatk9m4w6oPgnH0XuUzpHepPjF
a+b5M+I5u2odAeEl4MlbvbKuynhw8D437VI9Asicn+vxcSDXPwJOgLGvY9l3RcWyqr5oSiybxBVq
h/2v2KrCvBIXV/rJVR78eS3akNrjDCymP9xkgxH4r0N1tLy7klEuKuSNCXUCoClXoQixERoDc0Ux
+IfScRaWkY8u/Ht0RxdaeiU9cgaEWvMxIoEX9WnGk+pOThlz+455SHgmLt7Paq/LUyBNF5CyApUm
un4e3AwxvDhfDg/aCX+OIwQ6nGaf7aGaliTqkmsnBX8XN2bBk2ypvmfK68l9ON3f6fX6BJjrbAV8
QSoL/vC7kkWkAUUK8RZyE24entHrNSjsDy6hXkTGHFtFTt8/dnpbX1kYw/4hhUknp8DtSK6IHAqe
jcILNKZBbV0GHJ4F6kCEOMkpUEC8zuxy6RQW+vL2s5MU9Tml/jnkH0wx9Z975IHRxl6NwT7LjuWe
fNcqq2gBqOpMas/mxALjhJ3K3YWYgHRN3f9cvyVAE51jGLZJ65w5R/OUXkG5GrrYjkVSx9c81kA3
TjPHkTNZ4l4mfcXfiAIgrtdEuRXqdCGmWgYUoEXacJFQpBELp9I9ufhze4B1PdpbLrd/jW4eH7gF
rGsZZp2eP3hXYdBBXZ5kCHMDgU9YEIsbr4NvisXhEaFuuo4mOvGDomlwh9NxRqdHRhCZ5kJa+s+C
WAf1eJsaDMjYBcSi7IEWs+EaOCIEBEVqQsFKE89sUvWmMx4JjV+zFbLRhc3NOKSs7SgVg1/weH5W
ONvwQlCKK778T8gy3O50ykIoSQSVae2h/mWWX4FxjXQna/4Ar8CcMqlqcdMU2Ln6xebLsszLxXg4
5z6UGz210qiXW1DD/QRS8ayxEng2wc83ji/L3W9lfXfXt+wflV6Xi6z57LNNkXK8iXzZBwnryl9R
Bef8vkdqPk3aenIZtGYMGoBLtPyaxJqp9Rz4jN9HGSfksgf8jXx8Bb6kH50BIzrtq7JXxhb4PHyj
LWCb19vXBGQzEZOiIPDZwZ0WVHXWiVdcLj1IwUuTTL52QH/PUdW1xrxlktWIEcGN+kLc0HdjAurQ
oZOJSMgSPlREIKf0tdCg2U3QZsMSIg/RwX68z+FxGCGTC2hGmjRKMMN9ctvYNB9KZ8J3OoaVB/BK
Hx6md5PO6lXVVqJzW4ZHl1wbJygjrZcRn+Otz5YtG2Vq/G/uj7sX5UWvzus+5BGr84Lef2QB6vJN
KGYolMcyJJvQJo2JuA97lX94uaji9JsGHs8FjNy+q1nEwfvzG5jzengxqb4h2XuR87q/Fnrrue5g
xHXZayp6RH0296P3Jx5gKorgPaSFZldtDdJCwDqYcBw8evsjPOl4nIHSqie+IHm0+HkubSgarLQ6
Hxl/mZpDYkpA10uxlx3MekmZOpgfvMiW0bOGAZIC2aWey1yodJasPe2wDsHY6oeunCBr0+AFq2Rz
paErM2eqBMTTjJa6k3pnP+3qmbv9L51ma7bJbqhoFA9fvCwIAbSIUf+9vQ/qunX+7XSOhVJjS5tS
CrH0CfWQcbpkNyj7vheXkiH9qY2BOpeiPP0jE4euELnlk+Jv/76PQ+o0uQkKKqUk+D9IkLa0K1/B
uK51Orr2CvVohjgTBbUs25noWVDhrBU40nlRYuPu3ci8lg4lN63R1B/eaTc6cv9YdL3PBulk6e/+
kBmsh20paUCEZpXckI7Wz9PmOGPMOCBWNaKTCi98YyWhF9siTQYY8tuI9JWKY010yj4Q1ojeo6+F
LEhbfGpKGjQhzuUQcokBcwkXjUTae7cJZbbeumfusW5z/2cbKoiQY6XxTtbBWO+74/ypRrS/GyTU
10GmRDOsnN7g5vNa/PfsxBjpWhMO/3BjIH8xjkWDaNMcDO/1m1LE1DNHzb5R3htRTqWWlbaB0QFY
ZPNEqAjrveTm2qoztTvSfv1KYEq+uydyKZAMuRYLy7jnVoW5AQGQw3WEPyVKZ5J12Y72lF1stYON
59+eaCtYOdrOM5MpXouCNyaopz5/AYboqDj5VaGHrP0T/S69Ecrwtz6FNkrPdQmZJKBH03tzD8aU
GxhQizG21aGIYCE1e9EnMbcLEoErayXRPphMRpif/bzu+/AFo7/ysRdoqWVNkoBZstS2bqVCamzY
qejPeBSNkAhsgcrT4g9+gBYybeWr0jkP1P4v8Pf+K1Bzqo9LcOiK6fwDxjgzcXne9gwppNbpPAUc
09Sbn+lF6mu2QvbSNydu0vr3ec5H9JQiueehbCvreswFy5qHKgYqDTBl/S4+5UdpctQXv5NWlCtZ
9DHq5q3N/Wd4gKp+sLKuOdY32s8oFLbZGR4OjRVTYTWTwRGXXrPw4/hg33DkTgdh3yCMphj1PMb/
H5DIqwMBfZK51pOqfja8aKbb7cXy+VXXy5tYD2JcbSrV3UaHHwMeXdPkgke2YkL05v9cTsem/Ltb
d15ANwna5h/TqJztecE2shGQWaWiJwXoxnt4/EaTXorXkLzGHUgSJtvCWMLSJD51vB9B67m5cuE8
jXtjRp1gSCqIplW8OIj1xPoq2v9SX1rXPu6TpOFik3DbbUQocG+dqUHqLeoq3X+Yi8ePfP2x40rD
zwHHFTMyfhjUhQfT6poeAshT4egm5GkLcNuMQTD3ANYS1PkxXi65+tsnjKWj4azXsxOZc285hHH6
9RVXAWsgSpAd6FZTPhhM3ouBkimwc75p5yOF8VSGNmGmnI04cGHH70Nvtdv1QRmq5DaiAj33USxI
44K0Y1tF4uQZI0iITTCVngMHtIOhQBKQfP3Vv+mbqXeq8iR3oY6oKu5ui2VqNeWlrhf2fKmpvuRI
ieJxnc25RIaQOJuv3AUkzV86qHW53AmOjlZsIWOnM8Z7gL96ExQeVS+NoSVw9QBJu5eZ71CCAtjg
0zaVncilSlT1/2BRNVXMYZiB0AXdt6F2f5TgNH8/taMlqmYSDM2JQxOuQVImk9OBHQZUvAH2pdI1
PjmsPGdCEeeI2tg4hYU9gQVQymxt7Z7RdO98hu7gliamFUpDWrF8L9WcgY+zeCewSKbzzJEHxOXQ
OltDRLGdU6tYxKujYNMbJ5RPNU8kInMvjaypiRu3tI6BaN6+r3WXVNqqH7mMPJl9nD+yfkHhBI1C
siRF3oWoo3fTyLVyDKDyugtGSHSgCp/DbToThw/5SeeqGD3cgCtafK2YB5RDPmAKnFUZAfV7fY2A
48MLFBGjoMsnzkwLiv39yeo+PhW8YKDGOlw6Z7vLI02oa4NmZCCLSiTmolMBZbdAKyIyO32ey5fW
ozmVybZdq2y6vgPnC7exa2IicyAE3Wkb+1K8Q16u/wfGElx4CUd7HWO8HMFnqP/iboMzzT+DCWkM
0s8IFDzhnD4fg+0KnSVqVeAzySEiFvA1LJfQWebK/YQ7sAvPB1jkLZOGgOu4cqUYPhZ8zcO3gmiA
OKb9dXu93jcvTUo2RSqCuGyfmLIgzCwGTWTYRX+GwknmHhetUUXZD/9gaNblc/FjUyXZpM/b8z6H
WD3JW7wLxpNWwz3ZGUu8/BaiiEdtDtUueji+7VE0jBClK6gOEiR1w+RTmlR96KcNs8zzMgKDa8bN
zB9Kdk0Uno2aF+BShrjreUe70M+upWgsw8PHg46kYU9Rdfqj/7qcQuhcMjHiGKKxcKnVKgaCCezH
cHr/v5tPwaDEaUUGMdPPZhYPXFfIuIb7bhrng7F+3QrCUCABz+xsuUxDsuZGrNyBrz7ui6g32lna
I6kb4q73YchHwXKqyvMvn9CeFxA1mdrP8A9VDiVY5YbOCcMvUJtpWQrivYEm+Niw9zn/EHRj5gVi
TmuGumOWN8zR/8eNEYxZKrAk/0VKgu+ndFo1be+aHarRONNDnELEJUmgEV+Ch9SN7b599tw0uE/9
UicFoPoJSbQUyV3+7qNQKzZ+wyZRMd7mKp4u9wouyc/on/Q5RgbMFtKnNhHVriuQYqPJEGv0eEiL
ovIIJRd6Gkv5LQeWxhrhobOvWqm65JW9jz1NOIlR+EhaKW6+ROM4CDS7ndWjM8pB6gNVABPgxN6t
AE61WKEBKWwOKgnNtHxbb6yKuqgEFw8Y9vs7TAfQv1nujHEi45NC0kkO/ni4sm4RxSt6wljOOih3
VLiFpN5Aj2CQjWAzHRErfohSwhM+C7ANGxZiWDVfjIWMw/ESoKBx4GAs9i9ID+GzRpDJ3duWg+Pa
AT5n27sBFKpqJh7JNoMicRQDRbPuK2kyXDNHb/1EUoYi9+QZDDwQ2S57O5ggwo8rlfVi4KCYoykt
+K70Zlm4+FJ5aDBGbCzkSXojZChviINI1DXy46J89Exbq8hrBu64rMKObha2xSO8sczth1TGVeO/
k8u7WEhuxfOPlQtdIpZo17iAhrwbQRVcuFijgx5Gh7J+hMH73g4btDMzioG+ggMZ1j3Snj6ArDmQ
wzQ7SD07LE6rfMn7O5yKBwGyKKV8VucNdIr53uKBaj7E+Zuzk17+3aBZ6F590Ag+/e1xKOz1g2r7
VnwQ8E2HD7O+3qS6Zx6MeScJr8RilZCRf0+ME1Geg2ndpm361Az82Xpgt/bnqrHNzuoQPW3VGwLQ
aBLRl/GwN+5YctDyptp12HaZuw40j8CCLvCOVcvghjJFdsLNBeQzwL/ThU60JLk7dPAPY32uy/R4
PjEhRnymc5mwb6AvHdKxa6yPZejYyMqR664HjA5rzci/TDv+K5oLVK//JxFtMcyKgRDkv0Dc9Xng
zFIyA4QIOY6QifdcfgMJnYfGKCqtQKpwo0JeGJxd4yx//2r6wVaOWU8SU/+t4W0jwN5jKemyz5m/
7G82QPjyrjrH0Zn+iDj5Zb+laPcGdgPp2+qoJgZaO0+kyHheOoonI68/yTRpxENUUean82aZITUI
UA+ev1iS4ir0vDnu8sSxE5e2aQCAMNgF/nMN+9zqOuZ31dPkOErMNVaq/tyC59sZ6m28o4zFEAln
MMwf7CTvXPnic93v9SSU25+l1dOyIen420iBA9Igw1MLAHPdWQXCrf89idfqdZNj0dbtc0UCVyG3
TIuKdNZp3U/s0559gV245Z1dZ09wh6w8O1DLpPOgJOfJuksHpaDWadzU4UQLjctQ/u4fMlMLE77d
X1tANToUyJKmoTtosLKy7A+9/zscnMgJlFciJM/UY8Pqzzphvs0f4dWmjtvfX8vGRhQCuN2m8RNo
VQB60iQjNLoLw8xz7SF/+UeRTjV+OiFItFa8+t4AWkGcJfCFPg6twbsNFhABlX+Xdcj5ZKCD8Ckn
Behq6Oqm5s5e/IfoG1Uexg1Oz/3alyFjCwWNQGSPV3Epy9huT7jXFw1UZAb6LTMPVyduBpmUfYKg
BIRKzxuZHh1KzPe0BMcLySUTF9v4V2XxOVigEyZR5PJtFGveEinGurm/kyZMZHgKKoo8olcsi0iI
YdHsYnLgPs8PYpYVAMVDpGN7RYl2eKxDUzohPCkAtaEqy216KdWXxmOdXwXJHDb26viHVFnBC0Mt
4A4JC22SboqYCocNMe1hsN4NMk+JVBFv3nH7SVlZMojOF7eW5Qz3BVkuI8woaVSIWKYGlrfCK+39
X28nGMH7ICOFVA/z+Woz+xH5YDTji9Sg2qVh3EZsbUqbmWEoXTKSjrUFCFQIMHyMrN91+7GzZrUY
gLF4fV4ghooI4vSj0vroAm9OCqPas9ISv8CdDSt2XgGx3UV3Rw4Hk218kvC0CrdZyuNnJUQpKpZp
uTU6xXMijSc4lj1lGV08IBpbyMAG3bejha+OXW8Ipx+w+pIdi5GtoTnkCZHihO+mfeUltynQ2N2Z
+ulyoMY2f63WR5znk2VQqaHRpbCIWdPUY3uPNrjlMmnJPiQNRuvk/Y9gb27xT+8GnyMH0lMhk7+O
JY6jQFqweoN20lc2Rak3E8IlxhOPgJcG3rDUpI0xtcClQW8zacBmOkT1MINmwrc28Fg/HdJuUgCI
3aE6SNlPWUrjjbga7HZUT5cQP8pHlOu5cvI3PnTEMQGlIEqENuIJ9Ivxw5kmepTMbNNZcobrqLJ4
lnHJwfs4uSgP4GLG/l0yFGxW10iYUsERVPRGprsNVi4f/WdOWzLBdP9NLszsDymEoDXeNvp1gmOV
0L2XzuWv4Ot/59p3eEzuuVQjKQ4gL+p9aXh2NQWqzi1BXEH/VEsZBIiwz5PGYKSI5kCaRYsjcoIR
2+q4gfmKIwld1PSqCqz/+N5DsQeNrsej+0oNT6QAlia95x9OjAoXES+Royr1qTjr6TxHisiTpDNn
GsvGyBmEouFw1GuVTcK03BGERPPftpobmapMH2axQEAQRbyAgveYdC/gR+ZrZiTwlzrkZF28kUmB
YAAlltGP9rHaDjQ/fHZBEBZSNwYImcPDQ/tqaQ+ewBQro60zVVJKIMkjekuNhEEN4WkNOEXakgQ8
7IjQaXn1+IDeA/Wo+D0PBJcMisq5hRMx7AI2LqBP1DrR6MZ5H2JDf7L+yNcLquTQOWDQn6mcxl0f
zMHgidmry57AubAee1qM/ztLQ58Zbu4iIZzhUrMO0AjH52jk/9iTlfuQgJ2gfsfU210GIrsFcc9t
P0sQ7uedXixTxwbSUT99pcq0dT2gzuBHKT8peU9RsSeIbPsY50moDxL21liSTkzvvD+SecH1hN5L
aETrMlDFYK78sYR4hJZJ3F9WxsWpy8bRUObo0htvP3GA8R9bo4YCTKEgn8QmiTeVBm8fSRRrqRpA
tn+rZUysAOmZCBtNyh2zus2QhWdaC90E1kO/5dHKj9R8G+q9eAqvUJ/tWXCS2cr8AkvrBb0TUSu9
ovWIz1chIX5i5CHo1TPixNuGf/skwS23yMEfpR8ySy8tlZv/VwjV6HkG8FYYBxcmNmfzO+eEdI3c
63Gor1t9Rks3e2xcAk+fGHGmIG/axjreA8WvBwDlrqrIe2s1PqbtnkaVeWABVrPK2c4rjDZt+c1k
cO91X4MqsD7DKahVbONeDBbP8/yssTa2haIJ1AqL7ttaTVPJ0+DLqAfIPILKO7rasr6Bcc/nDvZ1
YMTA5UQ3OFrF+VwBBsndp4b8sAWGcBESrRjLW7NxTScWhAzvUcJeHpXhDdHWZSVDcQagctV6RqWQ
V2WycvhAX30DWJxaQmDshqyKa+WxCx9rnOmB9fZR92YlgTmWfVdkPDBMO2+SuFa01z/+qBRZIhFz
gaOlh/8aOKRu5oeAq1fp2MwGbXXGdndt/HSa8UZ4ZapWgBVfsSr9BmvzQYl2/xJOeFQ8QA6I3YIo
ERTyoo+rMmbjz4dEL8AdjO/RUAj5QjmMHIoU8sPeJzL4oKrvGvPeF2ncWRDlmSvGJ2CNFw+kTxUo
PyT7ICwpZ63aZe0egNRdkPniNS+amFRllj4OLu6tYcoQTnwA13UqmFyaXB2v5daX5RYoUaF2hV6C
psMmoWDBwmTPT1H66TlZio+3i5lcC/I+X2I0KRkU6Kntjollm79SV8xLvYelzLQTJP/vNP9yr2Xn
bTRAGXWJKp0mtmkaH9fzQQx7AZqj2qLvhpKXblqxqYnScpM2phL8vKtt+AnqEi6/NlbFhGqER3r9
2+v/fE5cjVJLDgtZ6VzFqwLA+VgRdUUirJcBGucCFAqHUyLGilVsKruNPjeRSccKHvhEm7eqG0ZP
Su32qHVs9senF3X/ojZxiPI9hYeJjhP0+upvha3/8qZ+wQz8z8NH7bjPKQZxm+5LptHWbeLR4CXh
Tpplfr14/FKbR5wdcB8qVFAW46BeTes/xoG91GApA71Aqq/Fv1DyptlhYTNwLrF10lFVWTIV/zer
gFtlab6U7+Fxj2G+qVqY8Ahtti89OPrBC1HDeHMmJJDyWRsFU4MOIPkWDqF5zlIrpE/MLaMTgKog
Iptk1My9GYCzSoizD/PuxtxxwhraZXpfnD0pBDp+OX78kifaFSXKiZJ77PQODkgeKNPEtTUho2zi
s2BFFPaPfE+XrL3Q1SJ1AmxFXGNXdIfVp9MiGgchkyK7UZ8Amy2x+8fU0aA054qJ0fmX146fZsDE
fs6+W+1bjBFamZeE9NUU5fVkKG1rZ/k6Dt3npmpB4cycgCu761k8TKKFjJ9pIb1HNwiLuuNuE4jB
68P4lkWR2bFm3aju9dVe40i+aw40ThnRkID9S6OfrMnlQEc3uXUKpNnVZEO/iOFvaySq8CaJwc78
9+QJQXVv+6vVBcphucRfzHn9MWKsrKXOFpteqfaxnlUbY/TjdkL0eSZyg12hYGBuPJUuS2hoGpHV
wRhCkb2r1ZeG29nYK0ItpqSIRvG7zWfKg7l+a7a9hug9zSEWvYeIQkNS2OdcLbf1CmXh7khJXnIG
//mctbt4hFVvrLssQWqGWGVMgb/k79ppF/ee6668zV+A7rH1Vd4PdDT3L3Y+1d/COAftGfE5W1ZB
skXOJjvm6hl5rethuWw6WNsQR9eOJ7df9MIjgUQF+sxjN7w4Rq/OXGOh0kQR029Mzw2R7wDX0UWH
wLks6KzQojsRrRk+FO30eeCYJPDsgAnUVh85U1vbRElanGSLPJPs1uP2Q5j/p60VSd8xqseSvbT3
Qk2o7UH0FoYc7IiQEE0sAtf7nKn+n4qj9hV2C5AgFh5fvdV+OjCxCTxcicvHv0Ib8Sddk+gY7eqH
SIPyslOYMp69FRzbi0Oyh0XR/EwhKj+dNADWBtL/1TQHgORcyuDA7WwpmH/jj9NWQNBkSHQ7T09r
ZPBJHxMlliJM6IohLKSy3Gzz0Bf5x4F2ytRQXi0KlruWHG1BBkUElTWm4vYnSbfo82zEBwvfw8/H
3GqJlyttAFeoTO9yYv2a0EKAu0Q5eip9kmuIN/KNnDknjhlif5rS9r1LJQ1s7ng1rvpZFi+Jxp9S
VUKsjHZSwAK6Tw3sMuSH79NB/jXhvrvIw48QJjkfnJ2t7buoReWY+vaFBSI2rXS09tIjDWNTNsJ/
qSvGPDfjZEKye1vayOv2yrrVSpCX5yD7XT/4fKNM8aEaIs0eB84qw6sz4w8PvqI1d6H6AOvNH4//
U4nJdbZdW+LIzceyyhh6rBiInhQXKaSUDc7MRZhJhinuG23qbi0x6bxZfHih62PH7FIs8bJmUtCZ
rQOHdDsKm2oBlCqGjw4B8pBpXPLiX80msB8lyRSj2gn8u52yd8+pMkrShyC6dMqT8K7V9y6xz2tE
24jeuQ35mmGIxOfM6bpN1CD3LCXijEUdN0fAVKOi8gjsDe4qXSxASPA+iZO7sCebl+k/V9k+d6Zt
IDv2icfmKVF0ZFfoGskmgKCw05jAWBObMiYvVUdtXZKL//EROVkd9dF2a+aq/bmmfxa/enCN1sVm
KT7wtP+oUT9RVQdcrjnQSbg/0ZFlX7JjUfwwvgn6VlJOLnF2BH2wtBgQx76DX99cWA+MuXgNBP0Y
TGbSPKCh4VgRwltn2bPrgJ70urZguy/gUct1SioOLXyOfJqKAc4LaGiMxdqnHkDkt/dUe5FmpsDP
3lYtGCSibaL2p9o94EOsk39HLSut0C3jGq1eSiiJcYkQIYX+9MLrmGULD8A1PLSTLMvoomXEoJ8M
6YttN10h8YPsfvwPwzd3O+BAO9kKWcBbcgB8LwHL+S+6EO32hdl0RRGnTDuZg4R21yttNFKascqr
bNlSaggoqJ2WkuSIRVn8f3kAn81rZ7OanG5oiDEW8EClRToRnJejUyTiDtd1GlJ4C0tbK5W6GZYa
3mWbqzePDAFUZKWeDQtPOSArwcbDEreCgjEXLPRh7c16hJrCorqREyH7PNO9AHgMH9fqiayQR+aI
O2ZnaQLTxv+x7koqgvmI6FRubsKdJRWbq3TiRo7+j7lOhnv7cu5YBRHjGjVDiXTwC9jr8bXDmbG7
YlCP5WqBb+9NT8/C84UK4NEuUmYfUFZoX0H81o3ke2B+LYBbSMILWNMUOLhZvjtRNp8XRcKeFV58
KjqiMPeWUWXMCyu0mmnQDWFBe+kAVaBMXQ9LLspRnY633FgtxcZ7lvtgj9oGUrfpbIa+Q+iEpEhc
k5Y0YEI4cKGaWmpM5vCssFq8/ExIJtQghoLPlILuZYaiKufzmunlF6DnyNbKxcyriVQGuYdR0KLo
1vzt5QfoG/K550kTyhip1T8kdDbI0yt7ZYRZ9OSSS1MJRSejwOXZdG0cWVKZpZGweWKakZMWoMWQ
FxR/kwKc/QtEAFgERZpvzCH03f5GOb5iePR1tHQGFD7jznId58xaaF4vxZeapsADtPq1hGHg9c3K
sP4dtxEh5w5r22WRsHstxJDNoYCB4x4qxsrMwgATlIC3Y8rryuXzayDIAT2bWlzR6vPwVhC/d97a
/PaI0sICiNp3SK/T025zOUVqd+KLkDAWBNfYFFJnzF5pvvynQLsOqlcNA0q02Kh3OixN85QLcQI+
YeB99cODf3h5JagQfvSV+47c5uDPtQErJWscztstYRJc+D4iB+X7CW4Ne+ZDJDZ43HcBFpXvft67
JpSjYzLTF1IWowE68xBGa03hixC5i8xUGw5TQyPP8hhZDdhCXRrcbOQAsO8hMx/MI3KWxIciytTn
tsz3SzUyC06jGLiTRmFUpZqbeAKmU5Rrjt50/jsm6M+bogX+ta2Yo2UtKRP+3A01A2jhUt89PJmC
5oiT0dJiAnudNhuGO/dIjV8+zzvrlbjsUguBwCZYlvhbZryK9DjsSE6vO64Jz5nSa+TCWbjIyjbU
B8CCkWs+lhpFIIcx5EeOrkLOvCtLW4WqQjUME6ZPCvq2QsR8WkssBzphubofl/NO3S0kIjYwTMHc
TIA6WftIZT3bIT/TZPDmVpsHEQslu3I+2ETlMkA/5qq7czrXPkBVEN+zrEGWyJdKQ10VES5iJ1b+
2PUWsvSyFr+XaXNvB3+1zTlpAejLKTKWHV0DjqsgxPCJre7tSJldmhG6CtrF1/x4jvkNRiG6M9FV
HMxZJdw440gxw8oNj+xihO0cH9TfKws/2DiUpXuqCv1eNwLSt/jDWkiRXDeqGjR2hT6YK/bavEbW
TJqCsoIonXvgAP56bexGMrUMI0JojF5atMYoEmPgi2nYJBy3Dgub62TL7TxwpiVAkeElt0hYCkSC
ROqk2ag5085fiB9gpz9xtq5PQhMqhMnvRviJxkOFbjdyPHOo0kBcEv68wYJ19KggEXmxnk1Nva1v
E5MrizJv++d68wAq3Ym81hW2SdIHQpaNa050qDi9hg3jLfaLrUDp4Hk+979f6pPhh1kIdqC93pd1
k6J5MJIoG62UAFxF62ElG67sTf/BwXHhtg2nkKuIc9ZUxvWk3YbXgEvP7L6kjVPW8zeI5A0vSZ2f
s6Zyopps3JMhbp8tT8TxEFRbhhM0XzADJopYrGyHIBGlYTtjkvVfnwMnfPL8mwHdMxq6fK/dNXMp
oqFHBpQdokX5s4qiGKdn7KDLmV6qTQwE961tTTgaPsBfTbeslvrf+6PyDGThybywVfWs7yS1IKuQ
7MBkBkD35BbdRnaD8a6901M/GJ4+9Ewo4tQbYVGaAlG6y+RvKMg4gtJQee1jsLRvga2fBEyffx6R
AP+J1lTngcwa/mKgzzL/kl1XmShxMbnxhJDeBKi7xABLfoao8OTa6sKeKgU8iMM3O2raC8JK8AgW
3j3OasJL2mBtVuvX7c9isd94god8jhPYkMWinJBRwHnPOXrZacMoWyPlbFOSC6nOJd+oyZS5CQAs
QjEO0eVktPAnVeSwzG+FeoW20YpduTGkNlTW8FTqBQTrfs8bHqESbWxKZlHSmDCe8z/VHwbmZ1KC
TTHuFczZG1GEpC1FoNtJ9TBLclTBivE3VoL8XE8gKtTMFEABF+JGxwZEGHxiWsVTaGllNPKQDSRO
nBwG9DHguo2bPuyGvfIvHZRcyZ0mGSBAQNk8liPxcWVzLdV14qS4XomK+GnMzyjkKoBiM0N2aJZK
CR1FrtIqOzDfFEUY04MSFW6/nfcUFwjZUEZlPHRvcelDIlcvoyL2nRL0yhQzh+XI7pXaXvL7Gz41
fgYxiSApx2z2iZyrw7xMbGlRlu67B5pCT89+hNd9P+O2f4vzhPahx2l422CcPABvWWHX5b94bWcb
AC1Yj/RSZDASaO1nyGpkFd/UjkYIwNSVpL15p5z136owW7Uz4ZIpmDWNTZQbONsnnt0TItqT2Jo+
ak8aWmIjSzAp72zzhs1Kt9RM23vXy8gdjBpvTl62M0K3WUjl6v9WXGnSkcF6m20OXlaX2Co4xXc0
czfpyxxwPrWdsDbw5BNa5XRZfD2rptoM1VYR4rNCqF4MjcxeydJiVOmxz9a6C77Gm++1uxzzsLf4
9QH9NOh0DQ1UI87TP+wqQl7IAcP1B7ZBzviwZQTO9jdD84C39QYdq66fn2tNeLcn41o4ole0Wryz
IEybGGR+NEFmSQo0GQEhBbyUW7AKhKnIbs4c1eY458MRI+SxU0OShGGhPApmXXLYKtulgYiTwSDK
Snu4XFXEa+A/vZcj3wub5wvmCKhmV/12MvTGCXQnL0r0zbLL9bwo5w8Eldi9E5JSacAvnE7krA6C
+UwZmhz3w2qblcHkKHYE8YH8py9pgzqCZ8oBAlIpkag+9pzISaV00VE+wg7P/WVVg2HF1Cw6jq9q
65aFhMYRt2HipYxK3zUEz/DRBcy4Y7FHN7vj4M2BaWYjMJWmZIQ6BX63SdHWCl9kvjaaA9e8WUKn
FImE/O2lpGfHvgqnAlK4nJqyN7rxoaxgafRYDt4Vwq+Ei4tnyndUNnetHtujT6B9tqhEYr4cNKDY
P1wOQrz55GkaADBnT/c+GLN3J8AeUa1f+IjHOwcXFjg7EEwAA3xtW9uqh4+rHID9HcTeXa1q2t48
Us6/yr1RzA1FBypPyKc2jGbjgDyRONBURS2zk88zxmi60N+I+j6t+KIkPyqPaTvRJErq1WQCj8eo
biYaIrh05T8pMZ+L3jzYZgcHjfol7yC3NVFFw7bxOFbcujK7vFvGkvZNY5QXrCct6zN5Fi6HdS/H
T2vijAllac1WOHZDMAxH9PpNzDnqvcyk+4hiFHDh73Y/E3Fdx8+3RIFPumgw1AeiNJ1BvhQ99yGK
SbhM1NG/dcLrnUFSmjslm/HS0k+06ZOpdoTXHgUcnlmzIeeomzv6WsAwVp+Q3GyioSAlo3/6OTc8
NMBu/8zjdK/M3eSfK6QLyUneEZrzhMaKwXzhRf3D+1mCwbDRru0NPfkJ4iMUvWpDnCxSIvrzt2tx
dTO2U16p+KE/vkTyxvjLzb3sJOY5nxZBYlEQ0hWemoeUf5yX/7rAnf/G3Eii14g9k7opmgGT0h/m
c7IRGfjtj1VVG5us2JZCLGTSIuNNnu9pRVCpdFa294IGrujm0XQXDBJlQck8ld0pR16Hhym1qwJ2
A3RDA4CdmlYbwstGwfPYMkaJ1sHPh/8aebPrGj7TU1Eay4rgUr8DAwD4b5jMdwBmwz/VWLN9G+vb
dlBU/D2H2tdupUf3CIBiYYh1uYwfyLxvfC4Ap3/uPuAkY887uGPrK6umdIXwPex4RewhdRht4c7Z
k5ypLQYWrTQ7ABkgZARBuTJfPWzKZpXOUuN1y5rm61eQBuWviTLzcdOrIJMvn82mEkQyL3vp3xMd
iW2cgeig4ZqHsX0zj6dQPyVjm4lGGpXJdF5RCraMSR4WCBStNQl0LNvEzbxy9lhC6ZWzdOjMpyMt
YTtZJ28yYvTFpxSmTNnY1YmIw8D55bluPiKMn2kuRALBCCzdJNw1CqgeZk94TFK2sI3fW/mX0P+s
vU2bZpmnE8pq3Tteh+vejRjHWoSdVEsnzdE02K4kJt+cnC8Av49OdoJF/sDNXAu8eRI8kgD5O0rN
Dbdwwxd//GLnVL7+SEcRLQb4JEFdtmZ+fcWhZ6vKVvuGJYQSD8zFV0Ez3IBvbOCC/+Rt8aUNIrOQ
KIFF4np62prfLmGG5+EqQbqrgEieDjJbsURb4Nuc0vu4FnAtdOU9oa8crTAZjL+WnzyRdKneU8/L
ueDnBtfWedUaQ4h72/F4rIespE8nD9MN451ymGektkhmyYA0Ab4ByM6eYxJGlU73qfH/zLQYIvMr
8jhXQBruFKw/kFJSgFl6b8cE3VSqEMPIJl+galJo21m0qGjh4NYnnsl5tBb2+ePPhVfQRuUAz2T8
71i2k5wtS5HWq3wJDTIVMwEYrPKagl5P/0AAGBeMUgo94fBkvCbBN6I9TXuE+LbRh+DhlB24guzG
tW4uok0y4UyJ/8hQ8lGlVFG1bTMOf/lY0HHyaB9nFzA7mLFEJMR11SPZ3g0/gUzgnRUMi98U7A3G
ycaLy5MBxYK0tGmJqrxOj6sxdtwQYGNipOBZ81RnEnEiZyXivm/C3FNp+uIgTS15qxp/B+mzo8Le
zeiludyXhx6duDGqgLwtnTvjB2r6NiXUlVZ+/ccK5UCDn3yKgWv1HJccAnDlrtf5xiclaPGAKh3I
yPhaVWKDQRuJHLRQWRKILwLh5Y7TSJOn8dMaHhBhLGxKJpI3XPQQky5dmH49M+kVICufaQyhcZcR
nvisIIYdzF49k520G586rOQmSFh0ekuT/o3QL+Zv2ZSYOIMCLXqp1JtNJPRHGo0MpypIi4jFzR1T
qbRFp3P5iz3x+WlCxzI/IUqJjMPjYwMjYEQR8kPdBfSvcaDyOd6ZEeRR4E935pDPep1sI/PNQfua
3MpYY9ZvzriIhY0MYF912KfEBLralpolDS2f1UZume2fjdJ52osqvorV3VwOOWTKqtx8OZUfx/OM
ZWjDBxNzA33TJaQjhi8YOmI/qpeHO4CtpjXJppNVw57JKF4R1mGLl+xx9+s7EfDGWeX951e70KXX
xgQ1ES76dUdjVwhG9jDQRnx9B94UF588Pc4mRz7wMfocbz1CJeT7+eX8PBjgrR94HtTXpG7fMf0h
hILXnmIoAIymFb2niZi96XSC4mHxsWu9G1B5PqQyX+g2h55gcFEyvBQ1CeEGrl67d3nYXkWfdKCD
/RvhYWlM90oORejpGVOkJ7gxhjhLXFmcieu/0la06G/g3ICF5bZEi2h3MT1Kl1/DmCj6I7PpsOe3
x3EUzaopwI/YtvPURo1vaBcVBYj7LpJTCvF3h3QWGXpFT8nV+4eXQF1hZtOz6lXXYnCG5FPEsW7Y
Veu6RZZ0IoieFqh0yu035lr0/wX4wfbch/radyfaGa46zwowDw0LrnZiMJiji7c9Bf0DNNQaT1PU
9R3HNuqhDdVmlUjTPaB1Sa802DCR5lrIMQT0/FTUOmwBAC+MewCx9CwC90cJQKpvwFcxnpq9gm/F
wkGvD5HN3/RQXkCkjE2jCn1k7sqOqwjzsVBPQzFtAsbovKHwQj6yRgTec28CNKa08nwnMy2jjPHn
pYxdwRLHpdSx/zrDUeZ987FdRZxoqr+nG3Uv5GmSLaI2qReV7nzS1J5mMh4NNYBxUxu6qQU1uLi3
sutI43uedU+nWRVu45GtG3IDem1L3/NPD+nK/7kYAlVg2mUBNwTwFQbevbKHs6qCJcRtvHvJhBVj
y2p57pFOBXjP/b41DVVExj1Z9V0ol5i/QnXPWDn5l0Bvp/evI4v5IowAjWc0Q49uDVt5B7o5NoMb
Yqhr4dlOYVn8ewK7rFAV77hD5RFbYa4wpXC/9rWwDXN2CHgXUYURp5ZtJw481sGRDogAWTP0bhW8
fjWoz+IVh3q1Iz87cgvVJl0hTVETz8Tiser9KkrLaTN84FKfSaYG5jkrKMP5527SwXiG7tAt7T4s
Fd3+rjqD5GRLHNRXnyZbDKcS3Yi0o/JM5XWcOcjtCOhFdZiUlgdYzYtaEbbi+oHgyEhmdXWZCVbO
VX5OEntOQRd77drJogTC8mkqspL4318CLBncXmkDqvCiNfWhKYqS433SJ1q/79lQl/t7fiDEm+VI
XdQjTVz366KdeVtPvHDLx+v2x9LWhGD/LbMVOp81dvpDn8NL6/1i55ZMjMPM+wNvah863bw8e2gW
wdkgiXfbeajkW45XHVTC1jgA+P0i9SNFiMcKuz6U+6SLGOwUq7pWGNPUFYNdmmGCfZUpdrtxmPkF
dOgUTSsWp8qEmTtvrysw/dsc7IPOdUDpcr31c9tJSI7h49618Y6CxEX/5LzIT+r0eyH6D4nXeo1e
7AbFH6drG9cbYHK4FvXbBsRfBNRz1NNDOduhcY0KD8GZ98wXtJv7bzuNj+orK5oW1c7YaxtV8sZE
PLXM7UaOjtzj87aiU3D7YzeSrnbISjcCbEUJx7Ujy60sTGLxEF8b2DK6qFSAJx2B3MpCYyhTPEfI
pRZfScq6fC8+VHd9yajdM/+nIn1efIB8PcY1Jlr+MhjDvJ8yCpOCq18zCB5BAUsoF6WnHdE4lSrZ
B9ZR8W3sRakgjeDbYko5/dId7zYpZnW+m++wy6KjbYp8YT1CfTCeeYoZKjkSl4r9oP5FT1CfDoJ7
p87zZrcaIjNsdz81U2XQJgzZMmIvewa2cs3McFcknUMaSVGRPEA8PmzDoBXjo+qfePH7tZ9J6es4
f9QfMv/yX+IWiFX8Np7t7rYLOXAzMGcOdLhldYy0BnYxnOh/16D4ilDzS6WIexbd1fHWAyS8XvZj
yWgy+Kjv5rH1ChpsSdvwLiygYtcM6CMcokOD2b8J5n/wn84KbotG1epS5iMHLS4s4sBXmbpmZwdU
yy6I+E1Ge/IO1R4RSC0kfIeHb5CuMWAsnJ885+czYSmTuXZYYRbD2eLXBo/jqMIi0gv7zrhPQPJ5
76C7KtXQ+46ECp0uTjwjCmIk+Nu1cMmNEgoqKBijTRZxzBoyd9DgSeoBhcQXOwW+7LjCVuCPGGJ3
Mq9pTu2E3bdsv46cnyuFkeLMd1h6XYXQgzB+f6D20lQ8PhE4RwSSpVEEiDRWagZKdL+tGbL/uz74
tXZU/AYrhZxLYb486WNpvS0ije1GtdUzipGSiYCbKP5jKrsMZAmk8EsymCBR3aKZCAmx7sdljLYC
wHRPktTZ5hYENR65NFzIGY509rccP1gUI/M8+A6EJnI9vMUVg657eChc8LbDiFO0RGktw2VUqtLU
eNIT3Lk4uWxM7ASL6QN9RV6JvBC+beVPexoDv36dkb5Kh83/+cYndKHNr8A2PvAjWXODhZJ1YYXA
pSS7TXE8gwGPveuyQmBIa4tSZGp6+WezwxdY3WfhuEc7QzOVcncrTGLoAOnSZmfpCJyodlrbmC87
7e1AlAvZg61KTweXM8zRtjLF2ufX5IvyDoB0NdOQcGRfzC79n2zDFGTsgB08C+RoOr2XkMCtcxBt
8AYlelhuxPdtojohEMkgcu7qq6J6nRL8VWVWdOlE8Rr6P6tspKtIWR39ky4BwGVQqBU2VCsvz1kL
TIWqII06+QQPmeLCTEtYoRT01WRMXrxZsNPmNERigGhqu0I95PE6X328s09rvAhvO7fiXKtI/ixm
ZrO0+OyQpB/m5wGXb+hVjhMLqdg/ZlZu+hYBu1aLNJ8rljO/oUFCc4h1MxhYnc4LTdSK1GrH/SW5
tUgfD1ku02BlFiEXwGqHQJFJAk4TtOO6VvvRccgFEHmHb5JMeiYroPQKlK80Jn2QLaYR7/f8fmyZ
bn+G4bLTVEpejzctnPuvG74bY0cwo5FiuPZDAoa8gP1lmOIalyHNUS+LlcAU1KCTs76yZa5y4f58
3nm9Wc+DJ24KQK0iykYNsxPLuAuMPAYsSwAsU+aqqut0ae1nYhuGDmdG1C4LSrDSJqA8zHvXy/3W
mpSmALwDOer5W3EDBvMqjYdGdcsIcI9xpOG41QfIsJLUGO6/KxdmcyJzDgDMUA4qshNVfcBoQxYg
z+Z1fRvZjTSzVEanTKyzyeXCNBvjnkP27uuIUcPrucLE7KYRQ5Y4+ZvpW18Muk2ZLddmruaP78RQ
rde51a2ZhkvJm52mFUu+JqXx4lb6uGvnVl6sU+P6NXzC/DK2og9DMFbb0PlUc2ROCGcroCFHkkta
tq4HQW/Qu1sJanBN1nv+EKBFOLSBvUEY2Vv7dwKPV8RcqW7ZdsxJ6nVqYwqqF50hea3B1T8qS0UM
d0VkfsjDNJMDqRJI2cA2GtehpcJU8WWx45ZP3ZmJq60nLqxW4+QpOeFoqXIriN4wm0zx3dlOsY8P
4pqPxnatpmG5+HqPFHRlJJPm4WBVOhX4PZFYrUbbFJQ7MDT8pgGIXciCCvScEZ3aagZqAlaKAxMZ
Zl575MsacbiriYvmqFVsHXSRg5b18KQxMKxkDw8XhyTeTM8A9qU81Xr9pTXhlXf/JktWqFSn6R0h
hGUU4j2HSKv/IqgZ6f6F0V/+QvTwJ3AYU9tEq4voMVA1K4QXMFrm6uQcMbahnPOYlNAQu3t6CiWk
RjTn1GOA3DxC5cVpiNhHSotccHjNjrOUMBbDfdrVARw/uXTvBr3uuVh5zPDdXIs3les0VhsobcNa
AyI/cumq3Y36He2Z7I2Nq5uxKXrW8HD8K/5aI24MLpCIm6YHQWxwJ65p+ZEO6vkry8BkpMv7FxLZ
71zkeiXQTUdMDbZ8LqStqC3mIOWs9FqfqCg4niWIrCXcSD70LOlunwRYuFO0TtnrDa57hn/J8UJx
arEq6CaFIJt00AqhQAGJxmzpODDCdtrNS6p6SpwsgIejpZNPOspw12AXa7c3QA4jt6jJxcWkJhc2
iG1qcjinS9uDivuQQUV/Bu8U1EJV76LP2YFrDTPmfu7euM6mMU0azw/wnwy9t5Eb2gJnJuZAOpes
DsIzCOl5t3kutaI7NhqNF2t/9gZpyA3VXPcb8lnixZ5UdvQvtFl14az9Wrsmgk2w/ce12d4q7AGR
PkE4Ah5PRDsXSJ6sqt8RKO+MsiWGv3S2+tuULP6JvBfpyauO0hYeqpCTkTZFgvu3bHhjrfnTbJ1m
cyCLHHutPAzJ4dQJ4/UEbXWydAt5+/BMlOQtFp2xNeOsOixYhEV3QFTQ7U2fKXQBB6lcLw+Ll4/A
FTFGUF0yJZ+6dMOoVmQ4EUoEvtFUg45G8hWBQnbVzPZLLAzJ1uZSwt4lTsmua1HAIhsoxL4hutF5
vIrdQrwL/NEu6yekcYVhgAFNL1YPjAc/6HdRvi87PWj681v5nCZZlq8C9e0rh4XycBbdBHy1SU/7
T/he+KkqmrSMXtKSyFu7/zCivAjtI85ar1CRF34FCDfXe6re5tYhCjdbVNSLsce+u+nWqGv3I6Wj
+mVsC0XCBEaTgcKD88wYgtOP/v3qcPFVkADKdALfy4c9ZGobaZ/orUdpw89E9qNX72a3OxAO+3/Q
0Yc2iSh3fgyLqVO+UgS+06Wx6S1Jm+nt9vHxYm1xuP3A54OPUcPrNaHPpDGEEnbIMxh/cae2eSJj
3FnPvbZLDXA8EhgiM3u5ItJiF9BYJz143yUD+LmeajLR3mvo0IMz7R0pqWe8mHaETfrPkxCa1Lrq
ItO77XGpOUKxPddDjSwNsPp1sXJ1MIYYffMbn8gx2249MD8DnE/eeRqB7xc/dgAkI0g1r85yQmts
as2MMjB8Y3D0Qa8gktACUkYwGS0cS2j3tEkcVqv3jZdwlMLECeU2LVs2lxVnBeTZWYLIDNZJdYbA
sEmAO3jnwQ1fesst8XS1SjUMuuPLAZLn3Dbz9rulvfJWGOacAbG3drgmmlgXJCzqL5O0DGVuTUwv
K9cmU2ib2m2uIjFyR3VffVeg677o4jriqwMMuqxfG6of4sr23iUcB4fY3JkMo9t2Oo4DjDHQCaUl
Zpo49dU3NK4vO1ATITEEnnDgexPaQ9r3Hkm+wAumWnmOhH9tcNZB4rhPnDgNM+BLcxzuXbXCc6Py
BwoVIOhomjRIEGaWt6Cdn5ES0G9wzEdGI0VXBXqINGnDhk6fqTKdt4/IRtIomMzme1S5DZT5dAxM
TBh1TknqIXt5VX+BWkemSEmN2HfvPpNN3/E4Z84lePlSsJu5wUt1G4UgIbQAFp1HohKRNJo35MaN
lZvSLtGJfwo/OGf6WA4iDy9SCpsH+xnOZpUR2TbJv/1hNtp78Pp4LRJsRWEpgFX3pRsmcZtigqgc
iXs8/hy5Gc2HxPXP1IqDDLTSyVfJ2MoQqbcpwZnkLyBRUM0XwN9mwlke2vZ7RquYJHtiUYxuG5Fk
SBjoWopZE8/5daNT5yeSZIXNc2fWKPzQOUivV51Qlw5YqPsYDHASi32THaqhUh4+HFnI22TXs+uA
B5tpulScNhlw9RgJtFAC/JyniqCKZHRVcxwCV9U7TcNkgzbcRIef2xDzc42Ck8WJPigGlVFnEGXt
6kk5GH0dRmHOaIRkG5weGApQnRke1Ch0y3vxbNCJR25wxUmkmXlY1b9GjJ3x1OF9A6XAEJeOo6XA
Cx2KYs4IF0Ft10OhNBPYkeKBYm7SZshy3W7kysYjJok+YQMr27p+K9OZaY68uJXM6OlmhBdYzP4C
PmAkrEQGAWfaESPEgsaCGoh87ggdPL4BS7rL5j3W8+KY4UdzmkZKm6cqVwZOSuIGO60/FdzNXtGY
1mKMfzf8gp3E9k4bFwaHV/MDFVQ+HLUMAcv+ZqNdwMYU5Vpu+zJ/yBai6keEHWTR8SavntYNCsDE
WVFjt7IFw4NuMFvtnVDoh53xJkFySUdPRnEhEckbiEdDgsSZDmDyoJgiXeYkweX6Z63kczRMzeCp
0gQSbxV2cPmOsfXmsWfzEYqewAQkGNQfVxcFkBmLarEA7yR1lockfGP7FGWS1erzZ30IPuSsrhDk
ficToNvGQslIvk1yEFRRLKpoMXlTuZ6xULBNvkndOBQROBNGqtwc8YfZbO14t4KZh6jUGYcv3k+y
qqENRWY3tAjlJ9uZkG9TvRxj8J7ec/5iaAxE1L1JzkxPvOC62E85yXlcVIO+K6ahsst+WMqDW0y8
tfP1J4rakxXoOce0P13A12PPN2ECEku8xAhRiCQSrue7sNdM62D5JLwExNIknnGCZiehyJ1HZgsZ
+cQTKAz0dU12RHiYfIfcGv8ecJ70bYjEIwIA2pCi6po+fzaqR1ah60SJuSXeFIE4JKD4RieCtjT6
ADCropEpx4JxMlAj0fnXXC9uonivXdIamcMxq85ngRB8QnNAYYQD9yMacn7XyMFOAOPndzMp9way
YqAf7uHT0gJNS5o9lpath2SwiXEz+fEplwYhcbxL/gy9ddBxoP1CXJ59HAvXF6NWEuG/78NQnL8+
9DRmSRU/daB7KSMj+mPXqz0EFUZutxpkrTVNFYc41WAV3W7DByzc60OPBC837kXAF08a0wex7oIe
Z+UXKNF9SawMiiXHwxRjgLGwPL87UJ5pqj8dFfBU3vuUaj11gVezOAOZbcxANnjXFafu5/bcK9ui
FUjP4650rfWPax5DTjL9puhyKdu9LwhjfguBUDAgUiaC8dRbSRDjVx5KX0dCOCKzfzM9GxdAS/QK
0sC/Jnq5jN2/LN4ZB9IzeI/gvcrz7JDElVNxfTTuK3ZU42RacAxc48+u6lswHW4KAb1q6L+nc+MV
Ra43QGl+RPR9ffUqlW9G9I5mQcEW20e9bItiQIr9KvY1rBGECeTp6B7R7j6KbYKeSGOsLR2wFo5N
sS7xh4uw5Hf2AQw0z/4G6inEOfsrxWSgp0/ss2vaTGsfkVTZYwfmy2PkWuoiVQXENdUvKvTOdroQ
3GFCuEWifV+NVbADwtprHjk8fAEHonnYM2mCngwKI6q7gx+ZIJth8yurk3ILiC/9uLuvEbKecccE
gmAoRv5ugFWQxvx9X/wSfti1i2/neDHyNpKUsWq4md+WDqdIOh2+/pZhA1BinwK9szdmuUv2Ga1k
6WgifPlqV87lweuE49X2WEeyRuPUw5SDWJie5D0hSmai4YakQBQnJuLU70Eei2tBW8NJwza3d7H0
Z/qZtpGQOLGEI20w+c/HLZ5TvD/U11qA7f7UafeiTkkIOIY62dtFUa9WOi9AB32X4yDzNLakgNON
rItzFn0rlbftC29FC0ZBst6LBSHu0ff1LV0EMUMpKz3yy99/vQutwz/1mBz/f+cx0c8P3lhy92Kv
DLGTou6L0SAXfYPlxp7q2tyceDla9feoIvpLaZEdZ0mD73OtB4cHOAub3HnpzrpwihjLD+hcWuyP
p5v3wpZy+eCJrGtDKULwoY3UI/REdfG80jJoA6UiVEd2f2pQ4WOBP79C2kkG8DTpHkpyTRYIkzpu
Gh1AWLY2Xn8v0kx2F5g9GIK6/5T5sf7DZ51kHCWFbpq4bOSO4tW+jG6wvhThPBkvMJMhvp07Uaxw
YSlDIMniLIPQGcT7DcSuUjiDCcLt9WOigPawwZ6oPz/N+qblW9npOVx2SXyheBD2rqDqLqdPodIs
Vu4pfd/qUkH1IAOgboBUtIOBueB9Ma89HUaTj36Lc90tm5VsUuTf3sYbqgwkpBHHpiuQ7wwkK57B
U3hqqzUR8pvriZMClsd6sN7jMEDVZmp+cETdrb+GrjzIX9BKaj0vWZFsw64pRvfKOLJwFhfzrQyQ
Bani0MgEI1cZQCBOknA6A4GBjuwv+0JzA4gwEQwQCv9O+dqi8pGOAbV+vRHhWJT7Nn0ADRwcP9NU
FFHqbpI8gS5K1jD1m1/vT/ywCk0WggPRzAwE8TXj1PRsFr1p+shNx3WpNvMthAkARTMd3VGmmrUn
AuhP3h3VdIGTGaTTFLAS1GR7f1Yd+Nntfzn5b+1SGcsvQdvLKeGGm53FXFuLvPH8Eu8oZL51joz/
bwxcjwd5pKnT6W+meXOpjqdWSv+tfSlt4qsdl/lIm4RmLPu5Z4USht47v+eMiVRP2d1wMVKh+YWm
dhK5WeB4S+UyQM/7qwkmK+BD4nNhDfO6AFDQQ+JImgWgQ37kiDrEGOCXoBI+VvCjRRcLPu6RLA1o
n34KOWqnG7fmBnZFMQkxNYnkYNuyKu+ZngQ6YHYfSdfuShfUnGXg61+NswtvTGE8yGtth6r4oOoT
Q+mzRgV1Yoz8pwKkKD3hht4C8X0nlZceZRHiOHmPW2VMtMImeVxcldahavj6pFpO3lN7839UCPR/
/QdzuiYksZB8HbycUtMd1xsMtNqW6Yjywb2Acitv+yW++tWz+KDtSZ6sOvul1M/Ebt/buWsI4ujE
gv80maqobCOPSNHFaRiP8dgIeCaSLun07U4NGfQPBUz1vgCWDvN1s/FXrwZfDoNv2vnwmGXSwRQj
v2Nesv2oo1BJsuDG9bLbn/MY55Av7GRuLLy62SBDTVoTrLkbPcmb4t+jqEtAFkvJXlIjgg8Z2SX2
50Mz/hnf6kutt8l/qIlonledo2VEs19dyfQfR15zEZP3AfVYbl12tbhmZ7xYXcNNH/c38jqeslDI
hX1f/MGMW1yRxDiXQpU4notKgif5LnzxNppgcvZcxD0aq0DqvDZDxTeoptnYcIAT5d8zk7NT6zov
3VbDi51jdh8Vhx6rOPdV+EpUxtmB7HWLhqnxQFQ6SCvaOtyX4Rc7Da7L1xEZlhJZr2+XQVHdiKvC
h/m2OfUAFUJzy7yyBOEuA/KAHiKl8BlzR5A1YDovECYjskMOMUSQoo8Wi8rhwANxgYhZbWz5jAnZ
kaPnrXVAwrcvt5DMXKfjZW3mZaG/5T6wxJiP4j09tR47Ioy0hAVZowECQkmgk9rIte7Vgm5FDF36
k7fSj+dBvqkttpJ8IJ3fGOaOF9VOqrhr5It8GUcJssdcz41yRKe1hi1YSiUXjhajOmNDIwSpyxiq
ttFxofWLTCIbpND3CCgTaZsFeObCC8cQorxDPGhq4r8kUfNiXrZrI/3UeSLC0ZPEoqs90xBb1Kx8
9R2C70jwImH+Vj5R3FtT7KJPpN5ndIQ7z2zPmTzlK0tlOmXNHlfPTrOXIg0tX5qDFvDpaSyOL90S
CCxWA3ymZunH5NPI2IO3AX9cL8FM+j5K9OQMfueEKyq3bvOuC0fEvXBaNfmXzTYGLxA3DdPaF3A8
Pb183sLTlR+PEC3kUO/q/+d3fU13KPrXXN7k5tqdnsmeL/eObZlmdAiXsagLER94Eh+6Jv4z7oPv
mopAw6RYmBDQyJwesDvgwydqQziMQZZvluNpJhqJeR8tQAklTwstevoQqsdkQqeUMt8w/yMINoun
BaKi3v87uzmFR5FMwjads/nKHtPI7EKgSl2OlySWOb7cus6lZ5NkHC0kovaVEO7TBO9EQRXFxW8j
ngkGxXHpTpWJ6PL48f48mSM7zmner9Hfz2+6eFk+RswLq1Lj+zmIM61VeT5PGbX8OVGKFIjlCly7
bIu9ppT7kc2ZNvRRkSQY0Q4+iCBep7UFWi+rbhLjP/hn2KLTmACvbPVZMkWKdu+2qjlu1NVS4cCr
BVttUGkf5zW1D90PTBb+TI/DksQfadHV0hSM3cB8HW87pinkJJD1If8euGv6cCTHfbkzBh2UndFY
9WLB6jo0UgoF60sR60h6qahIOi/k/Nfg8QFVyJJXJtTZcJE1AWAb+7r+PEtMsiC3bmHSf6mLNlRA
Y0Z0LkvRtwtxQK3y2E5PMazSgJRxSUqNu8kTGH9kW1TyjUlgXyN9j62wpY08CyAV55mIwfRtzpwV
OQzqKfTbylfhWTUM82aH49ewJojiDaJ14+wXTR7ITbrc5aszcoHRoO4Bklx6wVDiK9a0ZN+mYiTm
UAokMHeDbm6iGV6iFm3hZrCQ87ppJVHjXivbm7weakQZEW7gcYt50gs/QlI/IJVK4N/ZdF4DjFhK
dmvEFFLDLXhdfRcYaOkqSqDm6gR9eDSGmSpnpvuH5jUx/vjcNZYqc2YOCYwFCKBzKX8dTuhRj2fK
y9IPBFa3uWJfWqAfLwqBJ/3DcDVyE/ICKrJYBWrtDa4o1Zunpb+XQbr/2hvZgHf6KLU4VahMBQlH
OqATJJAtgRP8/tCcn8G6mcmvlJKPYzoKjqxBc7B60MHquT+KgvN3CFVlLK1vtCDEAjSy2LHiITrQ
LWoucTHYEQ7+2Sp1ImtyTftw5WQ6u2yvMoKv92GerYad2xG1Ki/J/FuQ/gs65aDbyZUd3L6sRC/f
k2lnVtG1Su4FN9Uce9ewfBsoT0ldT0X52yNgIYUtHTcmzoOj6x9CPuVzofyXxAeM7vWf4LvL1D/o
Zw4uFAWomKeT4WsS+jVWBe/2UuUPN466beKstnr3L9BTP6/dqavYNSOFhmvdmR+uQy3iDVw/+Pew
qK6zr1DowMJ7sncotCIBvMSWAgism0V3ouX50zQNPjybndknF3v9ZdMNItl3mPAOR1gQ4UwbwJx2
kBbn/biibfPHKZR9N+Jl65UdkcRm8MaoskKQ8ti1wWCqZ3hNLxRNFHUm+YOMWqRlOt6Bu0vDmq6L
eq4wSS2ev+/DIo2Ni1tmtswfvkV5LEEE9en1Vo1ozz1yKjAAeFQ2RQpguhcKcUM838ZVwpZfl1Bq
E3B3Osn2W+M4tOSRkJ97KN5HzaHCIfGf5vMo8agEQ4/hqqwu8I+KENF2kMn+/2vmEw2FQDK19O3n
DU9dv42A3mDCvHW3Kw4JZUnvjBo+s7fHWbl6KvPZjedG9Pqv0vC+2XTIKtEQCPTIgFH/2Ap4rY4Y
yWSvplfr4O5ojNOEfPafy5JBnBa+hvy2Bc1pnoQ4O6XdBXJ7keA9sBWBgX0fr8IvKO83jkdJCoX8
4lfeduh+GDb8X0dxwsVDrmaS97gTKdHm9NO7WVCBA7/gbnZa22mUormp8lgEJX2kdxTb7hi/nlSW
/M19molk6K5YzsIAebYyIOP8+fPcvyQpgWzMTXuEMHY43I1QZM5Gu7NFfkFKE2XBT3YBx0em90p9
cgjoVV/+7chdXEroRB6gj+4b+nBXUT9/w3UOxZT1kf2l2gwRQ2eZuwikDl8BU2GGl2bCFuXp0DNc
Fln9DKUKh+1vuHUb0DAecGeVPkes1cv+XIl77ia0sSTXwjwFYeHDBaM0UULZvzRdaBbTnKDxECJr
fx+QH0yJ1Q9REHy785rnIihq8oKslo0PKyCgMzGV7zuoZIept2hg7SXdUBup7G7smWoZ7SChsmCi
rUMt7TrUa3s8gSkIcbarNeKVlcPvcTZSoJBbRCA6As/YT6o3GJsh5Wit2T9gVf+etkq9spQEvqsN
XzfQ0Z/oHmYKvQo7bn65IkG7CogF6ruZuigaT7W0RBaVVl0MOpgyDMuCO1fsyHNfrEI5CRzMwbEm
YWGMK5FJhOadvE74qNDLaUKJ8/qkhGsPbYNW11c5xjWjboZTRcYdXceLnbH+2p6/qfkdQGcduDbS
Q31wL2lysz8ymlmHfn8ZMX/4N8sCDeqQj2y05lK3PdXsM6OR5t4JafNt2eEnLl/HBS4Dh1crjwEW
H9I55lZJZ8Ux+JdrCxpIOvFO4Z/XYTV4FY+oYfMYWNqPyemOE8+x2gTIxtUXN0LNmS3InUom7cN+
9k6eN4csZ/tHnUGfG9EtVvhfw02ihgqnBrbV4NxXLmAzapm8JaMDyzWEVz5fGQRjMpCz75jEgPCt
lytvc56WlqXkEUm88XZaTVT/IzSA4CjP8OHwvo0DtDWLCo6tQOtu1i7+LFsZJ1Ivvg+MTsGDZ5xE
OwiWfpd0JOQEqyjZ5aURz8qHyQUjFCrUWWzf6b0gGRi080E6HKYMOakSXiF8PSGpwBHNSqEJKDX4
zE6DvCn6mO0gXws/g++JKNCBXId3ZPW0/AhX/znkJDJ5kes24uHJwbYUFMQCER+5HzhoMspYKNnS
Kd/lnbImB4t8q7EvLqAXrQ+l1u4HcdWv5EZgdl0uCA4gseuxWbFeafUIIqGcU10nyaNoOW7121oc
sNVTi09f6aglZwDtFKJcXi2csF01qJIiEHrrfm9yjNeaNIQfUhSqQqxVWsRJ+23dpHoiNx9Cw6By
AsOJrz6hSwz7c5SsaYUfaP3gXk2q/+DpQLRFY3NaQ77R5TnmqWAEMZ5b7yz2LFa+wv1myS8dx+Cx
wSfLxdTWL+V5qxGStw+q52K7e7T9irWYTx43um3xVsQxAlzOhyATC+i6pxC1jXl6VlVLso2QwH2v
JLVVrAmVoBMqNwTK09qs1bzcWXCtP1Ve+He09qsJTONDy4D/iMIaHF1CEMWmuqbdAW9RmrIVjfxs
y5PwYpq8oxtAuO+RJE2xEryD/KP+BuWNE9L5jOC/IdUN8CHTB92SWanbHHAdL3uvHzaykmaZWdmO
ZpcWGzfecEaPNbG4OZvAA1yzKBBNBpYmUISsu+gwIUoanB0R5qrQQGZ/qhygPwwNwjkh9el8njkz
FlPm3zXmUzWexDudUKq6KulmJhoUU+7rFgvdZNV7Ude3rAc6f0m24To2UufHhcoNlSOxcqQqr2fi
TK0SHNJ7F6S2nzV5wWmk4gL4T0fydzHSMWnmoguyPqs706kU+crJPv25LRJL/PvaDl9dIb/XkuHs
GLjP33skJVDiiOa3ILR4n/ldjMNQxE7x+Ij6JQzjZstcEoU2sJNOTy7vojXoG+mcc/p5AJ35yKlj
wNOWe6g25kSMRcjTAr4Ism2OVtkXI01NlIhHXu98iY4BbrohoXlna7Kb9L9mLRjwpmYc+DY7EvEx
OH6TUNiNQn812bQGeDQ2cdCDcsLFW9W2Mdbv+CzGX5Hi00dGKU+/Y+Z2O4yDQm6YMtjXgN8KVg41
AAxowit2ma8GssY25d5WVEzItgmtvff42f1w3uMsJJpHOhZ+Kz39ci3o4dCTNt+G7vI22iK6+BSp
tKNZCJnDxSsYjop4f2vz8O93ViTPAY4LqcLCkO9iQ37jmpvFi4KiXeib+jZ2cjYtgLQRVT9NNZKb
Ogbj5gvrNuizSRihXu2CNeK1P5FJYCDNTe4iB+bz5lWIX+CTaFtvx7438TA7gHNOr9iTxSWJRI3H
MNP0vCVZPSxBh3TgQK021Zr4QxgHg75NUgOwpLnic/JTS6Zu0jifqh2sdYHjaxCW0lcYa5LWH5x8
YQh5zMm6OA4jEZcVdSWHlZx1ne4bN1LJomsFnCvxOvykB1LOPCpnCiJkI+B4CgQbIvZJw3JYlw0g
IG6BCpHHFYbvXOlHy6COshxuQsAtWz8Ixp9ayGKllnLcLuvbOE5+va7tll0+v84iSsPSHvuDGxe7
3Dug496hyLwkWUo21iLH3gMmjelrsQxd+lU8KR41GDOUur3tY8GIeQszH7vWSWOt0gkY/gy44Mcp
Vy271UPMU9ZQ4d5lBjIqi5Wc5HSSvTiRexolH+8ZKAWRqCw9RuhElHkwm6I6jFTodZKCeMnjAo41
1K6SmcYJaBncunNgk0c2dsox9WQp7n6YcSlUtv7ALZ39rnJnGEC6sKuPQRFM0anKIl6mEkmBFnT/
oOYdTk2ZocGpN/VOXn1NVzUgOu/vHh8amP2HioYIxmBp+XeO+s4XkjOi074AMwdAmQ83Xv1k15Di
RMWQrA7e3y0wNkhZJunvVEPXsjlMnbMc1XRGE64nrhwhNoG/wUdzU9mHGSvVPrXxvhH+W2K4or2t
bgl8feAQTIfNAUnYfz6zruetOiYFpK8gmSy5lYZFVdzvGvoQBUrI3vLwuzAw/7KpakQvG9mxR7l3
F6cMdEmh46BMfg3UXj5eOpdl4a9OCu/pxpt7KqKSoSfIKfkgNkxvo79j5tBu+EV3iIvQZBwAHGeT
VX9OkfgKZPZ4SCS9+Xc7YM5bQIsp3uBeMBhfqb3SwvvuRmi6TtBEgsdw0peYh577KboNpn7hkdo5
tJ2iEopbqxytzu5vNYtvx9t874Xb0q+NZ7lf51+fgbDQ4Q+1FA3IJ2XPLUfCHtKovoVBv71prEwn
iV+qngurgDccjulTqDst9xFh1BUy56Mn3URJNG867RaewucZYVR0Zdsuy8WZA0hueVL3a0znUE1i
hk4iknbke2j53WE67URByDGixkzZJboGBbSCfidmcublR31yyIePM5a+CN17a/E8vSogtl4JKT6g
zdhnr2/BEftcK9mb8yE5RIxK58oICu5kkBeyBlzCnRRj34z0D5S6JsSvWs7zmV8eTPZ/b+F2LlqM
I48nZ6RNtJhVXLF0x0HvTYaFKr9poqZ2eCGeBFLZjjyzZmY/ttt2skW1bShFXotEAzBBhva+2HjT
WY66q7SLedCD4NB//p+FuW546bhUMNYKRvo/SG0fyQtJ8oMchzBm5Dufq0CYmMQ1dyGUqmczrAKM
Wt7MUv9jcuV7mZaABefD5M1w3t21t3Scb90NtEgAxK880+3IjgH0jACdcFZHg7tFi5KVVHbR18+R
lG0yGugr6h27ZGtgrl4TWeJkKmGoxcHwRKxakIUQxhgBvr5ITHJTK2Y+Uf5csIxPQWIIyGQztxjc
V5/DQ1PPvQRLstr+qM4fqkVpAXVPlpnDJaq4wo4Hw01YBVd7/2W6FB+/n41XHGRL5YXORhiCqs0z
ibkWdPNG38Nk9BxNeGswQjFpYIXPGiFJBYZjEAlgXBhQVtnR+65j3uMGH0bkvAkDMGUWEHoARnVq
EqQGs7habL+fQAsTLg8AKAEdPXtR+DT80wffWm6CemRZ8Ho5k/m3wfnyzuS8FnLSJhadk1i1zKih
lWLkdTe7ym/XIblkb5P1+HVgL1U4aVhm2yg2KWz7V2I+dpjcP0VpDjaK/6f5f70gR31TeYi23M52
OoVCMQERJUtc/QvLLLG2MQ5LpXB/FVZvBQ8icUS/l/IUZ2ai34pRTdF4i8NcOPy0fyka+5xl66zW
pVTNSz+DJSbjq/HM3oT/5ELYYNuU3MG9xbm5Ng6cjs+zyxjbuFc7dRpcTwvXnYLi2AGAo4OjZLhr
8rl+J+nd3IDb6ubLTqITZTAT5H6hpmfmRmlODcOQWkkqngv/5DOyIzW9wmnNDWsFZi/LW7dZYroV
bJ/pHLPcCkCdcNQCc9E7R7hDVZ/NzKZSSC/N/qLEUv6rX/cysJ6wsrOmSrp7vfHQBcsnGvz2zHa3
eFfkTUt4GiNFHdYB53D0QN9vuGdI6rM29IdYysjpkLIhXZXFmgrbukk+31SR5DiQuJzkgp0+WZ1D
RNeywV1YMjIUUrM52ZRDDk2EA+CDG1OfOPpPTCeVBPmmVrFAZG+ImslKg8dF/F1JruYXH0XoIayk
MtGErseGJzAnYSaeS7TOpmmHTcCjWTWjebERuYuP9jsKIZo6ZLEX9kB44CqVk1ZQIsRL0FrOXcxg
X5zy2o3ah6efYlxoSUnM9kdMvyrieE0j7Q1zpVolLuiGcCbIwAqV8FxZXd93ZuFBR5MGZtybYklR
stdNaihJaPqJTuvf8KdwHGj0rS0ALJCQBWsCpeL1XpFnycXcc+M/JL0CS8gB+/ehuRnEWLj+VaIA
Hl4tHD7jfTAWEpclcXV6hvS4aMiUWmhSMuf1Tp01RBdUJRwXFhzWpVOR4MSjGsqtamOOZAVTL7C+
AKy9ElVyOm6RV4yNOV+qHL+YolhKSer752oD01bp5dksoLLg05/qcgHhSLPCnT9s4fMFKmp+U8FG
rGWfb0+1GefOkUb04QQn1H++p0CEcF3MnXm9PeTie0dqDc1fzRw5jUB5jav828gEe6N5XnqCUt++
18p/NhF5AFx+0aTbLcETIy14XiNwTjF5bS6k2sJsZasQmWwY6XySElHYlk7JG1plk/LPRCEVBoTq
MBkjnkpGjC+ot4tkM91fLtJ4a957ik6TZ6J7bLuLqoZmFwPRtCe8R0cU38ldCjxYtf2ALxVQ0bPS
BEUyh2giogfV4S4Vq0vOXTl6h0cSuEYTYgz1zZoHaccltQ8hiAn+GruIUDY8dEjDBsHpZ6us2VMZ
ALv6rox8bUEjAnIq56+SGIP5GnAJ7cR/bUMwWkkjg/nk/+cEB8Su5e11QGNCWk246pYkI2DrMuHB
qmDMxhPN0rmD4NqTJ1A07qiTbrjaCVoWERETpVLDiLzXQFFnZEYvoJN1BZSF87VYsTXJkJPcFN+Q
gQYl58U7VbIgwKqDdHwimpXSb5rL8VOa5nBjEPyXpoe9XHpxU1aS5qrEhIVBz1sYwLqICkNm8JT6
3nZi5Bt4ZWbe47u9MsBIqtb9bKewaGw7yx5yAKV5ozZNNqs9ku3KsK2qXdDIAbDXqLOl2K94VU73
Ro1lqQHQE3kVTif/X31S5qsMCO/EzPHNOVm5cwjG6wOdEDvjG5MlvBSogGcyTZQHNUP9YRxUXCV4
H0Keqg2db7XFpuO8HK/GDzuusowtNP3VTWGJ4qdFCMkcFC6s4aG8gvn6Q2KTEMFpBJmsTCSf0HKG
PefijiWgVmMEJDJudJ4Z47NYoF6k9aG0i6lDHXvRnW9UsqXgkhPFXEscJ2uTLLycSCNWz1Vckw6y
8t8WccoHt+XrF5hJ3BhuimwAoQhHL/MI9Qtwr+JTJgwqo+Q6aGbW/yyZSWrDhA70WT9rTpyYUjsR
l3l96rYYXRK0IyFlfyQuw6WgJylOFHN1I8w87vdxtPinwhEj+kQxIScTd35iH9vUxw0fESmcMsUD
nAGER9JtL8oKAKk3jWWXeFR5+36ZjVDVTxuoMNHXIjc6iK92TBS4YiTQIVnnXyus36CNcwgHKbEL
UbW5s26oubI2lm4fBcnbCJ588hqja3Gh2SwAXGONexFVFrvaVL9zZCq15vz9W4kWdAIgt4qZ3/It
pqrzYD/FUFJ2mirHuWkchF1aHSnfLt0OEoshMYN3wSbwIhOBJgsX0PFJ7xdgcP4tBW01U1JRKL3Q
MJ5MG1VGn9DH+Ha8cqTZhA4as+FOsKqwbqE5kEYWVRNabyw0xiXqclw6+5DfZknzzH6TF1mFkMjW
KnqsMSdt7u9RJd16RUwx8ut0XujMj6YthhmThV3VRieEJ5U2pPivovydtD5dpV9C55AFW8CcMs3c
w8F1G+D8O9yR30sbcIj8/lSk/RwuAKEfwZd4xDxwtWEWqt5coHMlWAz2OoxKOPkowq4iISrSmh1K
ESbVHI+7tYhlYhH4P70iY9Pdfd7dipFDs/dmZ1PojpadRmyUQx+YjaYiyyuDj2eanEaf0HLRgfv1
wKZU/pXt0NPQCdSrS5WABKQA5xg2l3IrOFEkKAryu1oFP4Tp70+fA/VqpHW8VSUd2Q9ooYs8UyE+
L7P9g//2iAzyKNVT19GElH6Mfe+aNkeBSEjF/r0gPQSgC7ACwanaXsoWJdOjwfkt14VAvvIyXu2o
nLc/7miOXfFggou/yTvojnO9Xc13+zzFRdiLzoeeTbOjAOEgQUZCLVUQrgO3mn+3ypBQ3I8uXfEq
JNaXhhQZlabfRQIAG78pDYF7MPVSPwd+6XXLpxNo+rG9mNkuD2HyzJVN0ufbEdMqccTqI/I5Lzmt
sjmctKcZTHRAXT7ezkR7IR4N89TWsqLHE2eda35kGqVMvlz/7BCh8jkCFPmMyZHQHV0EncqvFIMD
8jawoVdS7XPqyHCJcU3Q6jiJDVwS4sFtbTCPe/KRHvQ6lnUoqcDGgkpn5mOjk/QUtBgglZgb3FTM
WYKmeeijsLVC689dX2DLwrBDI59VrFjmIBMMsYWcI5QPKOmMW6EvxkO1fiIYvn5XhlstXCjE2/Ha
7m8MwRj1Og7nlNzno/cGUo8w0zxyzDXL7dosXOwLzKyJ9EOjVy4O1A/eC+/qy/njkXO+cH6gDe5C
RQCj/RA7dW+EZqIDVYyLsbZAqQltg9700l0ITW/i4NSvNp1YiAqsfz1CdEhJyH2bzHAZSqh5W2+G
Vxgh3aVlyyLIU5sZjS/fwnLq9agGb5RUPqRJ9n3XckZnDWX/B6NAglkMxAqKQRLVy15OiVgcRgpU
gHCEJCh/DuHEn6zF4y3kIP3AY4HtqWoGstJTmwAdgg10tgTTa8ZgdSVc4nNgnze2ny398SY4qqAH
4Je6Y1VcCp1R5zB/HhN3tai0bdk0xAhcX82cXmCIYkuOnJSTZpRL6wRv2qAPyc7n9Obdc1mPPmpK
gv7m+6r2tM+bdBpYBmQKJ7XlUAlzDB00LPk+3aByjhrZni2i9jKa811B16wrIUKWrSVlgHWsPfnC
0SOTisIf+ZyX5lQwoUMHqV7fPU7xaibRzfdP33naGKwREJxYFojPdcWcvPAO4KvOGHoLo90QEHm7
gy1G/SPeRMfIbvl1RklDu7eEieIU0+uD9yZ65H7dEw4DMEN69iiEfoNPvEFQvKwEoVtjHMjpoQPO
uq+GgxD8EpMVExXUomXFWo1F8C2pHOn1Iow05PVF4Djvtfx0ZsJlUwsiUB99F9htTPhut6GPH7Qz
IXyyG41iRV/0J+SMZnV8r2Z9DWqbPcZKlXkp9pdP14eFGLUbiinbuOLe+WaInUqWo3nCrN2XaZix
O29FxovJ5mTQN9/cU5nejxxoFlL9pmmewTHrmY6KwP80aSArPc5Kuo+hkV3BkCH/76OSF4nJOAOw
o8ibVP1ZJqFymwg5ylfXyJUmcol9x3MaF4vMjY60FZdq1Cj08ctgrlRgmmab6bjf5eck3HC+MhH4
tuX/jZC5qGlEAT7DywAkP4VWt2ijxcS98YBpjWF5e9EiYJ9d7P6LyqLXCVh2ia0vetUZ+pf5IVJO
W558BX9ErzASw98aztoFTGyxDOHZcUVhzrPs5KeKR8ToNG9gKvaQZBtwqk9gLEqfRxJubQ6tS0OB
Z4+/7daciGB61fexupYh7xOuM9DvIhEe11wP87EvR7XCRCGmi0eFFyQPUn3MJT29sJt6P6a2sUdI
eSMOWnFIExCq8YknfA9RV5BkmthgtNjMbbSgFhXAk1NeQn09wikK6N/afZKvX7Bei2nUFyuGU0Q8
qHfM4hn0CruCbyn3fiO9JDv77cM9k9Lu4mLWBlGaFhlMz2dJ7H2UhGkPNmm+kCBNHo84D+hU5fLq
jQqh/qVC2e16bUYTTLq4d6Er+sHZfG8UXgD36EZJu91nBaF2aKTbU4k9RGULrw9nqhbG53RmRuoA
n1k/zvZ4JoNx2/fgKJaR7QA+qOYh9z40Tg1MzHnIc5yw5/mF9JsHVlUKCQxDo9mG/WT/+F2yPFSD
JGl976dMe6dioCLf8unYW4uhVeb7anw83XTwzhX25rTsvWE0fFJ+KQZdkbUGdSqIVAfXoEUtCsuv
Zf+N/OorNw90WQAvOgAmn6zpTmWiuFhOkFp2mNVUsKha7V+WHmY3lCO6PFWW9yvrdUKZ6ipmyynk
VAJfHoEOh7ZGqOljc5sBIca6rjWOOUqiavE5wQV/F7UfbsGn/AwIudJe8iTVnxyCgvQaDKzxKYUW
S3/YVBFfSxKLQFq5Gty98qb5HmyQxjM6gGdYvRXrCcRmI0Iur5SHs2FdPHlWwYmsnfk80onxqbSE
hYsaIMAjcsl6z2gH5K8Vh7dyPJGNEHVQLlYYGZEsknkJ8+ViFIkhENXMirxYU0hgIEbxRME6CS0+
GtCQFTV+b6cLV7XaSFOaSYy92yEwk1Z693WYE2hgabwge6PoRw8KaevSOWulBJ/lnzOm6DPH4aDE
ErhBQc7vWxakqRbbVx8Wfja9vQGQ7pTj1E/tFCncdZglsOL3Dy2YHM9vr3GlA5bJLXb+SzOSFtuI
f8+gb5H58CznQ6NqJLaDilQedS68rzsUrRXX+UTwLEMWXGGvOlizTM5gipyXF0isC6rkYCpxB11n
83PDgP7WpG0CCJhmQqtieUNSbW1X1yEC9wb011wAuV7KvZr/eJapKZtYH9oJ/AtchXMqiUxsa/dK
u165N+SamwIthFd1sr5boc5AUMCRR9UY4A4jjYJqpV5wiu9LEzn1JCHRKhQYOttvBvS3omEVHizC
Jy1at+ZdO9pzex9b2EeWIA6JSaCFPUh1KvrvAA8MP/g7BgvYMUjo3sfcU8G48nep1lfGOP9TCorU
rHWU2aFCBsqkQDsW9a0B0fcvHOCAzSdYRGD+126ABdWzVJVVkO4902c0ep8jfgAT4D9Litd0CMub
y8yimwcUpn3aEFMQTqlc1FmnLxHUN9nJYnrgZXM2dDm4JPFRL81rVF+ewJfjWb+ZDyvPAqDlFhGl
G7KxA9MSIjj62+fK2Bds3qEH1Pt8VFxmVBHqJWupTuRNQPUUsy0wEVNaYw4tfijJkJjSDG746nLu
Fiias6u8RQxBe9X/1kiDKUwtVskgWDJukqgDvKESBbW5Kwqz6+WSyoM97mrE4UmOPCnIJareqCVI
l2tDBErOKcaVmnVNPsY9rU+kEZ2maM4MgTo7ntGdhLtMVREOBW/51EhseNTL+qHk2zxhZ/dB2z2B
h3yZEGhxljw+3W9kWvzH1+qy4SXYatmiNmU3y+Je97Y/tM3yTCL91/qADDuXRwWbJxh/YjY68Qsr
o6C0g3Nb6JW5uJBEQPxa3dZTZExo12znDdhSd5opjZ17Lx1AqA60rWK5lhmsEgggyMlff2pZods3
lBJ5PxlRUXJCCpX1v5wbua3iUlxoNCL8HqHOFW1KOoelwWOsEOJDc28711bsqyxSFjvwr22SxtfN
Y0Aq7xGBHzjHqopb6ma56uuvP3GqfW8tHErDdbrPU8ZxjpE3jNBcepzJ2119wdc8uPfwF3tr89ph
tlLwr4mBy8/kHynhq7tYFnKvLluoxO16Unf7S0YFdQk0f+rFJNG+Q5I8eUjxZzWsy9L9huz4TeUa
uRNwRvtCT8NchNT45E59FBxjKX5RxNsJGizXdjWi53S+2kqS8zkIXh2U8rScmc56MGrgNXtSvLev
YTgaKm5Ag3oi1TYw0BANby21Rk5JcMvn4yB7f2ZE+7vye8CSlrZR6VqczMLvppMbmQlCW0EGVs9G
BZDYDjqgrRDaY0XnbcxLwVzqT8F4JZLgud7nnbFEJDh+A+so7CvSEP8TEQjHI6VhPW/nn+jALVHb
QAEmVwQKzYyQTA4vLGsqjp8ZP6n+XVmar3z7NKYBwOebSnlvhvQtlf8yi9D3Iyyl9VyQUSnwIfuO
BqUyTSEE/IYCQ2sjuKeqwcjhWXpf9be7DXdfuD0Ez3U+92WU24PVaMlDwO7MJe4Mg19NN4Jta+hp
1W1/sx558pxgxPvlzIleUsbcE9QEraSGVzwA8Q7kFvN+hrhQjlccSVRpA1QnzCfuVK/7wYsp/b9z
g+XhKIQWYSJktSt2SPRhnT8qpyCwrd/7n7bb4R9f9QYF8atsthEBCSIlT9Hp/ekXE0IK9t/REt9+
pwe0xAqfkqMrqpcpvy7ba/E6oAVqBeDNJ4iCMVAZ0X4vB3a7/t0cHmb/LZDZwWB7I760PcETBce9
4k8+DNBqE7iBNQSl7z/x1m/t7UgCYH562cXs6CtKJjAAJg3zwzw/PeryOPUYyM8nNrLoYRFn/d+u
LhGcG34KjKrjPc+lKbJFFHKRSloL/Cg11DZRQ3aYfyI4oeCFneR9+ZtBwuqp8R8RpcMRueOyUdKB
ohxut32FmlUdwSIwIj9j9XIDNAhv5Hqb/lQMKj0XJ7XEDB9OApfPyyH6ofy1VIj0JGXka6j8mOs2
yaFP1oX7jxnE5d7k9CdU6wPdLqNpgwF/4WZjQHZ3jmCB6/grQPf+1S39YDgSLZ+UQF2U+Ksb1cBj
Bo97zImNkXcG1gOyZf2At7YueF7mGEev7iGsBt8Z23c1MoY7tUO0wncWy3wNsKxSpA4L01F+GaI0
Xpco9b6PLx89sMjqngL5i8jksYgpRTVsWszM86STaWcvhR9apRmS51Rq8XoTdqW44o6nHS3dSWHA
6Itd3EK5C98frAVdmFxX/uF9pAmBMD8p8Juaxy/e46/ItUe7HvUefhIIb+++Bqgmr7qJ8tFLg5oY
JGAzB+LLgtEDuLPAZCJdkh+NcBHXsDD8/X/a7sw469x152IrlEevVvBKpxTxLI+y9w7bZHgaBjjh
YdCuLDOb33wtAN/xvmnPxLPUr9ZxRtM8k56o5w0l8R9457+pCweDcsxFUjeLZpTbE7Bm7ppRSlUg
jZAIxn8D4JhOVefbFXWqpo5LSgL84cCUZsP4ntqfz5ckLyESrHLoxoAtAiCZB2+2Dqzmd5BwogEt
Xg+ZZ8PXZ4PnWw/msRrhqb+OMpl7xnp9GjGXjGrqBKc1MldKIDVTzl3RS4h7dfaE9nCPTNmG5A6M
cJEWvWwO9u98oVi4elE8IqOpxN+jJm3j48cpaxKyDsSYx+fMX8grY2UmGgX4NjxYbWkcoqt6HWti
jhnG+Bjx3edDG8Ybzj3SNOgF3w9zBpzA/BxxkZrnhMcTCzQRaa6YzhseGv0atOrhF/QzN6azBMs6
Hw2TQuZ+hzqsPm3o8nAJ5B7trDS/DlpqZ79c262Z6Skf14g2jelzzquEXi3cChWzo72GVmmMHkG/
Fp47qrWROaGc8WvF0OLNuISzcrZH4tboYkl3kFj3FyrMvt8eTqNIXOq+LGDZ8EipUvf+cRDOoSE1
iHOnIkepnDafkJTHnZCLoHeKkF3sEcQZCOiQDh2IdLZjoewXHJnPDy1RwfVqWxp49VdtZf4tqdzJ
jA/gtEOQfUteKG9e3zK9vqMFPDcKhDn6Hpx/IP0pr7QEe2tC+h/ydQ59sVsxpQV6KsAveCzfg7ff
zySfIaQd8SCQrAQ/HV0z74VmgFKqTiSBSFHGLhABYxITE+unEOb1y3DWLG18SyO5UI0DtIg20DP6
jLHwDAl0ZIce5Vq2ce9i1IMbUxEunWhVCM/RcXJqR9J3e/nE2XAw25D5EWrRKxCfE/pXabK4ISFw
Ozj5cdVlC2eubmwQMEIuxBKKiRSl7XZFtwu3A9jTKL5YqVVsD9UdaxSXEe9vtIti2ILpMBkss/WY
QAcfe/f0jTw59sz2uhhlr3WNDIw5QeLG+iJJortTPkmLwdFRjirBCZCW1IKIHRkV6Q9QZ8bCGn2e
LiojRNkjlYSlrV3HcYJCeBkxPsOmnyUWVV8hQJTxI2/9fUS1heotSDUpL1ThS08j5e1znen2gfOu
L12slm53tXeX7h0BK0qwWhC5cdznku+bcT1fleHeQ1hBPTc1uuwzW0nylfqe/Id/5XhvGBuWQEGU
ZUyR2ALmTeOO4I/NAOuq2taZGvjOb4TjbUak0AfsJBGlEXYw65r8iVtvo+bkyWCeuaOMZdbZ1N+i
gbXZK7qB4cv0flvUGG1fAUc7NFoqxlq3KNn4JVO++q2Yd08U42b5LFSkXMv1swml5iOozC+FO1+H
u3cXrvkcAQDVG6Bq1CfyWneNhUy23D4GaM/nIKVNLYlIdQGfVigr5pEIgxIY2QTtpvYNzoIzcCK8
0ylmysZedvIW2CH0W9unx+5OXL3pSxqwf/WHfCT7sYHLvkdyTvNNZTVtfMOrDm/E5OEEL1is37/s
r0tp4Y/10eAsQJIxPJ5JpGAJJzDOa2VYrSbvnVgJPXxChbrjPqcpf9npj7f9diHcYw9co8+1XdSv
XYbpwXJ+B88vVGDYG5KILGuTAPdAGfAGosDhKSLUy0FnP1pxsMRDwFGaRVxok45XH5WMhdmy8vUx
yF8V8bLtFM5y+ltjL1fHeTIsOvSyPt/w0C7qVVAJVOJCZ0d5htNxoonYrRZZ3o7p4Vl31QpNoB9n
a8jWklmutr2mbJ7kjeMv+CadpNBt8XrP4VeCtoB2AqnSpnAFr1+1uQ4P6qjIjegawy88l5DWXcMx
oS7LMOionp9rvw/z99RDh7X5l0jQ4Y4BF6WRmkJpyj0hVBjKHBoUBwdqChOX2SIwOrD74dsvyfJE
FQ3r0ksj7NVjwtYo4UbKr7S74RTz3rtX05Tt52PvkQYnUFhvarpEgHPHOeDFol8abRghH9kJpluX
lO6IVXYxJj9zfOCmAN8tcMLgRtss4PD5FqdB7IhIWHFihnGmGL5ABhM3udMSr0giboxKyswTPktq
F6noQSukICqcq2PizXZudYacm/owUTyIoYl26F0m0JPoOaAl0u5SYGwUW3VkVXmDBN0jh4mq2BjG
MvLhr3bJleLNtdpuixNMA/t0tx+MX85d66DNpGfQF1/8GHhrPCHmO5gw9h1j/rTMDsEP0h6o/y/0
EshWQ8FrhdV0iZyyK3NszVumTk42z9JvFYDPbabwngMaiAJ7DaUD7Mx+P9lyoAPOFL3hs91eINAo
KQpt1rBvcrdwZclaOiUYf3nLz8CC15LrT6b23PW0SjCcmkR+EGHNUFglNePzDg4xZ6GyGDGRSkuQ
PD0PrJz4sU8mLCycbry1U0/QazxfZDsxycZRHHBpR1oIaUztuF3wgL5UJxOIlYjpWjWxE4nVuFlw
3EP6ESBxQ7mQWeSeWaY8j51wX1+uH4x01IxAqkVJQ4Jfw189flhczxRIip8hQg4LDDUFf3jmqSe4
MOmzJvi9leIWpjncgjtiaWaqTWfoikXFWnm5WjKzRHD4KUEVEgdBEMIueqppx8hsIvbLBDaAQwsb
jx9ZzJuXrrpkD3lo8AG9jmKtUCOgyLQI8B5HUI6qdgAazWH23aylu9ODLuyY2aoymzawca9vHmD7
AW8mxm2h5pgqnkxeX1Bx1akTj1GwuxCYP0uoSIbTVn5TII3Q+LCzabG584JM4vlR+7PHf3xB0I13
Fzkh/eYlNGPb/OixHN30wQax0d+it5EPm8BM2a1gMTKL9Jv067H9100w39A2hJgYFA+p6AsLzJmu
V731dHFkfptDTHKXOvMzo6Q1MM0i7BYHV57VOKMVbzZOdX1ECWuRWixfuFIQ/sD9y5FDb1XyMA+4
dNlG7BKDHuv4DFdXuSmvhbo/phEuuMGGGhC3AxjCA+8bLHd+4DcY/7NIMaAwsFa3t2DPj4Y/aL4A
hyaJgqAfTbF/mTJ4efB8bJnLd0nkQjbHHLbXN3WtsmbBSAbbUsS6j+IeGyM4AWpx7M5DHhJemfdf
jnuLBnaWc2I5wMQpaVcHUZZuR9i7GhTu6wlsKfPqaElr03mpt7+kZrqo2XQCx1nS8z1SitGm+hHC
NfpxLDnJ6h7GZZUpjiN6fV1w8XKpNa5dphcASqpYqKcikAQNyzAdsEsmCpXSDnMT28Mzg4aqY8wQ
dfvXa11nD2KQ2tseAH2Mud/sa8Cgu6Q/Tv7qep6o1TuB7V+ZnxBRHcHGt3GuvksppcRYM7dZyUnp
OBBAJ/+FFuOghb9iW6o0SfBZJJt/vim9YEZnpQZrSKy7JyAx0+sibqv7VyBrhoueFYNzhYt+lCBn
E5y3CVkl91lb2nC8V8G7eOXZL1TqlBndlssklnnt2EsNcEtO0012EPlDkjqJLgXfC8Z+yLnrKWPh
vi5vahp1A79bRNMVpTGn8593xy3/RO+FCHtGhdcj40E7rpSCzdmGlBAUGm7GZSU8PUk0ABdV7s6n
3w8C8xVr3QlRHUC/whEFkzZLlCVQqm/qHpG5jSTCTxjkyuLeEFJGb0/rGCD2Z+jsMga+trmZDHfU
LE7sbo2AbsdwL/Oo0InA/UWK3J5gqPNv9ai78yquZtp6ehaVVOWBC4hoNMtsgCnfNI1n7K/e8cit
0raY09uqfqZNCVeJW8tZcgKTxvfi4f9Tdfxj1wXtfRl71rKE1PDHo1tcesNzCsCAva/zr8mG/K5F
ypjObw/3mgCvKw1iDNW6VpdX6lvtPkJvn/dTeuAPuMyqGGyztdQW9PNphdepoM7SYT8xVTHbj0MJ
sE94ZME3/OdORT+Cn0zsNIFnBRZkFIuHPPSZAzfeci+3vH7SsNFNEBrUet+dJ7WBEOhmTI0rSqmv
i7U7sUfe9WRVCBog4utj8c5EWd9JjDHjMJGlLDrFoIKQmLjrsO4Cb/Tjzu+ktA2W1d91YHT5hv26
oscsnrYMXIv2VfL61DbzYkUpg9ub9b4Wb9S0WkfnZBhDRAxw3hc8eOmszIJ5iCjsfNLq1UuT0Wj6
j6S5A2Jb0JOM0EN5SD5RW1X/d+Hu8MPbEg/9MX7xRv+kCLBwviI0ewO7zrDu2b5TcpMGnFJK4ZS2
8vAKcFZ2L65yAJyRQMNTdjgyp+tpffR90mqUpc/COHJ2egCVSRgbDZw6PHvkcHxnWQW9DPvT6dk7
/1S6Qft2UmfxQj+Dvb2a+F9AhQDv0YtZDl/5tA59hlOefrShu2bmWDu+uzZzl9/fconcZePl00Q0
zp/4zqzQX5RHdWwinDwmJFB+Sng6atEZ01wPNd1VKAeMs2Sl3Rmp48yKKBxx3t8f0585H38LH5+u
wNduWho717eZH0GqAY+INkmBgpOEJdmPXfqmfZYY189h+wEHkPj6H/5GgdIDMFSQ5ZSdSOdIyNL7
wYypRfXyOs4bEF9UPsnDSF7uV3Zj2qGpci/MZKUfEALgS0Pv4yAlfMA+0ocuS1JKYgWnCkk3C4AQ
4c+4mI5gQvbYlhq8T2si235SFn8nQ3AT0L/FbjRE3D4XZNB0M0/xcNhnAAP/FWnaDTgjnjnc7WYa
ZCWR+BrnxdLYNgitWLUQPtVWMKsO5ptlaf3ci+QOG5eJXdxpA3NdLAaFTPYHcqyUTCA/MWQnAzEB
PDD70NF29esdmYBmhN8vChs0PjIVdYkLF6zQGa9FwC33p6dr73LMhBHQk1NyugOR5UD7k03NkegP
nR0B3AvHe9pSJdizhYrmscHM2hTY+kn0Qk5Q7hW9r3UgPsSljiKV8SXuvCgJcN/82yEHt1Iit/yI
tAffbp/yHuzcI82kmcc6jounx2fodxX0SNOvaIy5wJK4OMoZNgAVWxFNRJxBYMYnHMpj7wMwp+Bl
+2L9b66Fg/JTxKJ17U7B6T9ZkRwnrbRvsq+d7uCmsqUWsCZSuWGZwALh9/zLKY5lQNvJRvzMMUvt
tNVvhdJXmyZ2nfG+J+djR3a0TqS+zC+waJpH/r7cDWnbv+vUkYzcUQNALyD+f20ZD0A0nIx1NqGh
txgePn++5nYUQHfF8IIPgqJCXCujjcyk1l7i1CfS20XjU0ZznnOpmyT0US/JRCcUiJQJHikbZWN7
i+M/g/BpxsXueqWKYH1gjXFXJeIh+m9K6cLq6nmK503CCm9X1MhHC1HKKU2T7D7GhoKFgX6j5mwu
k95kNdqrdZXLdMUvWzxxmPA1S97wtCjBSxlB7FRn5mF4+I/T+Bi5H4i+cE6uOhH1bp/8lWsq2J76
KI/M2Dq/K9dub9cz4eBxO2qzhlXJpx37er9xMhGwa+V+3HITZdG3KU4pM1Y0SmQiDpeDEUp4/gfF
LWIxTMh/1wALtNHDD4n8F8KMSHNMwWXPtu/ZY5eAsnYji7QGrhmWsV8mqSZZ1Z4tpID7p4wkmGmy
M+5LOhu0EMd9eioR3hSzPP9KIuY5nk7c/uchu/YSVrUV4uFrOjrJXENUE77nUWuxUgInzKlI3km9
fRD/MB01CmLJvipsD38y7iQ1E3NMaJPnNuBwWt3ZcqpWih2X2eLSHXDWnWjbmcG7+K5TJ8/V1PUc
CZseHHqtjiM6opmXuaRRjZAL+L7ufNdiWvyt4A1akF7OmxFHmm2WXpEuw9XkGHXIfae+EkyWtMtu
EzJuVgLNOYOS/jiWO+8qU08EVkQDExK1K2TGzDCNuJ1fmEGcmCg6hwVqAdeCyxttQZgkWOuTHk83
taSFkPy1vdHHFBiKnTRqBjaNTK16VHPk9MParQV0yY+RHh5pb6d3K9ev9TCtOrjQg7+9L25NSvWf
jRyuIQqDGcP8ABgbcRE8HIlK0I+Wube9KnAIkgtnZzTU+zNMdnS+aqU7cSvANLOxwyP8iXOU0f3P
CY4NqfttC94jubaRUddvJMaCEyAwfiV47QmTyMcgHNQiEj0suAnJKWIj7neCIHrecXkgZyF30cI2
dm0xo9XBPviK6PEiwwlE2b9uf060VxDm820eJofT5i6Iwr8XnqXINz+iE47PGuOiQO6SxSx9Fbc2
o41Q+MztwgQz54vXC57e/e5RkGVeozSru8aXBTKH4lMFGRY0GQQxDujdXSOF2tObrVhXAwgifZr8
U/cUGdC6kUOYVWhZYhOXlSBxRr8toMJFv8ATqPre6DhMjlMGIKbD0L+YOC0/hu+qM1EdgUiVE66Q
s/dRoodbdO/22FxvL0BuPEvE0t4AvwTFTgf4X204ZanYGWS4C/J+NAe5QGRoOfPk6owKj27fP1Nl
l7sIw9yYnh81KeUoI8R1x0NiLP2Yjv+ZM1QPJpggSog4SyGt8HEbLdTCueBRILMTy7VVy38I/Et1
+5KI1y4dW+VbowalUrldGVQN3aDrhY443tGs5T0v/8fLEFTEuKStBbZOmCugGX0Vv+LWY5CNf1Ig
/GZT8UcMbzsCdSyt0FGQXd3VRTwFozlTap1EnQfLxLEUcHLsOBsrPlR0ynncSIY/63PSXi+FzK/7
75YM9K+hqxqmsBBWHCL3ojlS6pMLhlzmP1T3yWFPaOn7EJWJCeRwdHpShcdwX5Aedf7gf5wHNtTC
RyVoBMAnsVsi+ONVNdeTAvJKEygjnrW8yE6jOYeCI26kX5f2unqEAX+lx1DXjs2prI+hBz0cel6Z
E252TYJe/heqGgWmYw7ZwiErjgFafmRfK0xUJt1awirRb+ULmLfYBd/Fre7ipT0YocJMHDLZ6qrT
YbII1TLYHyV2yfRDqhuiTFUXKtlit1qycRWuu3AKPLX+6zJ2/0ZXdwHQurkU3v/yLygSyhZ4Maoo
71nhSv3V6pEJKaO8bopkfTfj6lh2YlFazI1uDcn5vgt1EhAklfg8paDsCI/32swtUesEB7eHS8NG
7C2HoI21YA1vmoLinEiaZ59XoF+5Qmr9gSyAgB94jrzdz/9K9UQr+1Ws4gfOW92X5qMdVMLZMLsG
SBwvYwxpImW872+25uAtDL/l4p8aATFzL+dlpJgVk8ezkpPoZwFgcExzRiwimESEEx62b6V/7Plh
XutIWRi8upIJtGOXrHpv59b7y2vLe9nF1WpPCKLFkQd98o0RvWQ7uK9ZcpA3N59IAkdMa5yzFBS9
ynzD/3MI2orgh+ksqXTtOJ9wXe1KfA6t/979hPi4pBCi5/79K0fVn2blkSjL6h332LQFcnAoKHOJ
zc8F3ltApxqAt5lOTaHNyF3l11EVEOVf0OLiXIe3T9bo7k+zZfXUhZfT3mt8vlL6oyQTr6zvIC9e
YWJpdGe9kxwKaw7i1VYu2iPs1BtTg1bMaQezMbFUgOd7LW/JRLdbF4r3rWTLoROIJpHsMNhI59PD
2woo1s21Om8VKAPaIkDesk2L69sRs+1e/qJJflp7dDBFq1pzMta3QAyZi5R44LKIFjgsX55DqEvV
/Yosxj9quabuzbVoEtLrypAI/szxvMV8Cbn28upA7AbwEwm2i6WO1z9wnRYvesvECe1325ha7zlc
gzgaczadLwvCxSTrmUEiraUd2zFxXLBCzNC8ig3spn4Bi/myUSdyEd3j3/NeU+Q1nSko+35YyIgB
I4FH0FiHx9F6z7KMcvTlL+Fq6ezOXlRGPd7a51FNYwoDB7AuQwlnU2No1fh9GjBDpanK+krWUFJu
PDY7iMWnAftOG5H/VpID1lTgDSzp/NfUD27U0uQ+SRBvP25d38C6qWsw3BYUvgam/9+rgawW0oAE
LOZdatcMJ1tClVFD3Bn/DjA10qAxh/yKC1xxKEc8dVEJL55jix1Ip7Z58iq8wEyDrFDt+EuCqIbQ
aqtDOxn/OmamSAuoJzJuFCqGI6GLvuBnBAS34X0pKFbQYs6MSA7YB8CO198wuoYfrs3eWtgY1nBV
o3XqufBktLenGVm7y5oPUuQlLJJPHXKe3+dnTMxJyCnL4t0H2tUTF8Qvk+VRKXN/gHDFdv+DKluS
//cCtIgBGQxSykbw4+9fD7O1MgL03YddNF+yN6gWKotmzNQuj7WTvtI2Cx9eOpshJbI7DPa7TjtQ
NnyAsfI/XMIXzWHWFL3KYo0oyHHbZ648d9jABZbhW6xQNZgFiLUwzauPKgNu3GcrfHviO2Lb/85C
6673AP2ibAGeGVf6X1Z8ieuWp5qru6PkEngpHWp2+oH4RyVnYJvuNAylohHrR/2gmeXHkAFQzPuC
lz0wWhfqaI4orlzBjydhtQKu7rjESwey1Df6GSq39QgNL5SwNTf4G1v8Dz96slaMIcn41RlYgv6k
HeX1h3nFGGKjUCYtwe6Fb5uJDuBoMpJUc5c82MogFEkNOcGvFzcMzVMNqYUWI5xGanPYoPsMC3WH
XITZWBaKl4wWR3bUkixtIu8UdvHvQ44qgZMUXUCEb3CixaVKFcTVGfwIEJnjZeL2YpNJMeYqq1fB
EESaqED96BxvgXubyAuEkB/ukEp9HuDarfAY+REcVlELhb3WP4mWzYYP+Uxwmv/Q51TvtptBi76F
e4tmIpB6RIggr1HLY1LAVWwyTWBMQL7CDRW8YvyJ6uCyBlDCmdyG66egM1l+Xk0tlfNLDk9GrEBc
kTRc8XeIJTzOnhE5HXMqHUKztY5xX0RZm+f/K3aoQjdEu3OClcT4ZLMNgI4+4ZPtACderAAZg0+H
qiEtmIrPjVc21w9WmS7IjzaWOZT/Sj+dd91wCmTTbm1tvd1OtwkcLi46O+d3ba9EW7B+TEaasqG+
egm4O6NEz/bXJaDBMMP9YJL3Tchu0o+DuPilEhHsuKKhnu4+efhp7kprNhzK+jdUi/bFvJwN7dQo
sdF/uINkZzq+7pIW4f//O1/WLmGd3Qa66ZKwWba1Z1PROJBoBAt2k8HJDV9ZtpXXzoDP6luN4QOj
qstbLM8AV3mcoaSF1165kd3PkA4aBECrs7ugasm58uuebLVKU00etcNmk9tVcoNZEOODigqYajpZ
dURXqrY4Yy977LcT8Vkr/y8V2qIZQLRtBjMbLPpcn3fVjt+E3ao7Oi6ilUzVJBLRDm5AkjCDqkaQ
3zYQ7bC/v7mPw0xWdG+hTdte4vtVAIXf8n2zc6PEvdeVNlUQlpglaATn9Va1EYEjKW10DWuYiIkY
KHotn1MfH4usNUAhzjzLVyMYGt0L4ouQ7PraxK6t/wbdt6nYlfuibo35CaBbUv0PKfY5g95SosQN
m1V+K/n8ZRKDNbyjoGAhirG/Kkjbe8NsESPAd8/muDmMOs1d50Jo/HoN06XEd7hrW0mQmU9THVLI
Brt7nzXXmjCw5VU8nsMLn/j1wagzEz7bYZp2yBTfjLV5EPvbPlh8CoMfVNYqe84WIWx1PwIj8dCk
r+zhxXXkVBbgZZAsrmc95GWvGWQ8zzlt2aKQw/4NkzBic73A4v9z7dyugsEyiG4XIeXtUUnLSFUB
7tycdYBx331x5rHrRIr7cS5jeCVmq14e3CITKhaR1RGu94n8coBhMRo7BwXku0q9rlyj8sOLqjWP
w9R8h+NqH6ff4NO/9P/Ey0Fa2Nx4rRLyCT6EjfwhtKvCPIcqD25CvLxV3JtbhH5vMFHie/5yRajh
ay6NuodxWukHHtwL+KKl7fxExAPctRmaaHbBy26kihXSVwbxVIfyPG9LzhAYXaD/eat7NhACz3u2
0O5yD+MtU6FM5KQYhHy0doWt6kPUbYeCUOIT+Et39/dtyYRwmd7c+Kt67IjtbwOIq+GwaD3aurZH
DWPmgXvKtI4Cw9r05p6jsvyCrVwIHKOBo5YZ2p5/0zqEViTbkKipKCtSbIoj1MSNlJSMfGoZ5Hv7
VkS+bvHUGIMD3qsax5JrFLOsWlpYX0ANy641uT0Anx/pdVDVRnWVE7TNJuhbGfA1NWYJunzpUlBY
C6ZhEEzSdm+sZe2k7So2UaGIiCXUUAvO+01ClYVy3KpX0/M6nFEyZXTmB3P6AHGpoRpD+o6nry12
jrEah5abx3ftnuSUJuSeWEwdV7x+og4qI0YNRca4zHLzOSMOzRkjZwyZkbzZfN3Va3TJtM/NLBXl
0jzDwmsnAWvHbwa9kknPZQTfzkFjYxifXsbk6nR3Qknq10o5GuOgCfx0/rLeR0KVHxpfuvBzG4Lm
tupUXyHiRdwlBbNPqBmDb5BoKL/Mc219FdI3pfK30DlXTl4pz5KdfOAQWpCAbulfeMTI+ZKekT2f
4FOzJoYWnRl5Mp14LV3lSiqthAN8JedMoDMI6RIkwNh8fJkjXmf4wnU8QK5xsdz4Lta+790toCgH
gtwR92mITmN6F1PAGnF1Ifij6YKs7hQNWdu/Qv/EDypEy7ZGFDQkIHi9Sq7zoM/hMnndUy9FQ936
LfL5sD7a0c2mScDvJ4uuBdHzoC/C7Jupbuze1k14Onep6O6MSxJcMToyfd4PAjwhyc7dpFC5LmpH
UkiUzAS1D+c/uXNsBI6r1yG3h9ZQfsV9QCz53GoY01MCyP3FLrMNMH559bQ7OKNJdmcYM0JSF6Kv
/FqbjgEQAX10EOTPsulGY/mkH7T7AUZHN0TTyYi0p5lZRSNXOLJO+emc1Tm9XjZZ+4LhOr5lsvWa
XfsC3BUaOjjl7glOx3LhjtTgARLzcPk1ZfSMd3WOXod8559cgPOBFumc4TXMd7hCezChj2wxQs+7
6KX5oFTqw2HNUPCqTsEqkONf5sY3Rf2Q5HIwO+lO5jhsRESZ/8D/pc9gpCem0gmPU3JHOcTxCGH3
ph0qN2dVzMUmgeRiyAPkhSu9YxMVUYeRnDxoSdt8GLQPf15xMkylJDWZcqutsZ0P5KS2/1UlOCrZ
zaKZkUozdSWfLKatLlhVkH6i8465E1IY/diRRVqhPfdMW9joP1fdKgmj8BgxogQjXX7k1j7XLXNe
8ddXB/az3v4KlsarnR8Hnp+fadeSzTu/rxQqPLQL5s2fIBBiG0QJg+Hb9XJ24W8YAKAhPBULjLQ0
+Y5btuxz5jK+l6+u6uTGkRAw6GYusO7j75WB+HD0QCElk+dpY211yKbyeJHGuyjy/f7Qjh9btNKG
JLJ2b2Ihy7cnMNzGUHa3v6B51AOLgKSXNH67wgj5TK0B5P7sYCKuLF52uVJhW696gy0dxY4wfnrc
99934ueMF8nKJjbBpXD9nzcu4PgyzrNWdV0kIi8rNPujNtdkrRRLyx/ewy64VqNgOqmuo+OMDnXM
xGojT9gc0fVjuajztKpvkWSwtGb3QqOBmncdtpKsNZi9ZPN3rSLOBu/5Or7RjJLUjlC/mW/LmmIg
2ZsuCMiVBYgDCcHRLn4yXiSrha974R7DcbdqzlO82Xmg8pG22C7sX/pDz/l2oMklnWZMmDyTSJVP
EWypXAZXaSWH+QupPJlCra1JfUojsrj48wv2waysSA99rA7qZBB63s6m0GFb9FH6y9Ja/LPmhlpc
KyeYbwpoItaq6HLFLnHC8bAoOHTuJrYKoCrAs3/X03XAg5gUHPIfihJt7akOgYXDYZX1g+lh2D66
RkDbSAqnJdgdE3yakZymI0l6p/miiBv86CzZc5gBaF7HOI2dDy2f2fQUXr6ATvbzHlIBHXLTRZ/g
9bgFCaBi/30VvcxoaXhNCcCdtEE/+k2RJSv06Akr6WUa7kjv+QaHxeuxgcX0ER8988ud4qknjYf1
5wqxmRiFAN9g8MGLOdRgQKtBZqaGza2KRCicDcLogfryp73vt8MMlBkZ93+OHAmrIQHCh1ewS/rL
XdC0e31s5bjqM+eILvDxrPrDmndm9P/4+TkBr4+Nt+jB9EO7RFdSRqsleV+UY/QD/AW8DQyVDNdp
T8EAGoIh4COkrNwIigF64Xj26aNswCIta5Fmh3INakKOp6HJcyO137VFhElAK76zsq63kxtNiggL
D29vhCLZheuxqjjgi7ligw/hL7w2pWqo+HDe4sTCG9HpDSER8SgDHoY8y56MRnIt4TFn7mxF2Bjn
bPR3zTXxiQXqW49BJQw/g5xkuzwD2PH1N5STIyusdozBk0SGrYcGEyLE8yUzG2o4JW2mZnz1bTbl
B+lKV90ep8totdwA2Jn+2BWsg+dTIlrQD5RmPQt9K0EUkY+zy6GdMXJtvDhPVnpGajTxyUsUqAGI
A/7EyfkMQm3L8Mkcrvl/8fQCrsjsREWbkxM8SUdl9LXRJEVyD/3Ij53Zay1PwntrjnkqcK69ufIV
YkMWOtpGC5KKRualAKOa79Ab1BJ/TKte8YSfr1g7GTcHZJH2S8V6qr6Uyb0TDDyhytAM94XGxfp2
+jTxmTqGA1L/cOIDiENzSpE7kOIpKw3Oi0fm0nsQCco4VMecw9xUFBnoJPioWsKOhtpidunObHHM
ir6urSWeHXML/wbp7/2rIHjl8DIQV2VnjrOftfBnsgAP43Fim55z+U/WdRK04pghXxR88sJU+7cL
qiHwA8foNVPFYUUNXWw49iOJKBWD8gcN2xmN7YxTTsNRN5sGXFYkuXjuGjYYRCaRfsu4Oulxwub1
KIPdpn5T1x439cafkeqeutyyTnJnM/NnmWQfE2qXxoMi4kKRr93UUOp01uJMuzpbyogK5Nwv1v/J
RSv0STiaXkOaBCdHjhLc3Ukp8qmz7ck1aFaro3lU9mVYAgTOgDd9hFF708HUbKOGwYsY+XwZ0WNC
pNX1b/4q4az98CRSB9C7CalBy5C0dU9iz6VaT7icJnTqUooLNGaq4Rk9XevuJvOAkk7vyB0a0d0i
HfBhMBtPo1A8zlML3NacRWggqvLRDr/7CXe68J1LEzHT56DNoTHvUzgZuK6wKkKyPD8C/NG4XWj+
pw+O4E7T/BNjrG2wcjK2eLlPqUd++DZ1hcMJbOaQc5+O5U4qOebaYtU72hg5M0WPDjsXHKVjpVxg
mDoShcfA3OMl1cU3qCGSlqz95saY3hofJxjd2DKAYqGbJSmatWYXfXO0AUGNUZw/RAPPtHpOInI5
6BDhLem+B3cqvJyZb31XRrxo6QKZd2BuFpviIdr9jUoBFpHaw2PH3o3N5FCSqf3lhbsmklSDmgrf
lYJmus6GW3XbFqlPD3FmuPplQSk3/PXWOLn0tqw3iRYlCau60Ssy9zJah01CowNDCJe4En3RiIFr
6zaF3Y8C7nhPTaHLF4S04mJ0X0XxEo+cOs5xvDgnKTMGeW+V/k5xKFslPWm3SWK4ED8vwLSBRNQp
mnHFTsY8zjxcg9gJ9wxNPWqMRVaha8lNP/QirfkAEVOy3vmLKb6uLfi1eeSjXJ7RK+9ZfeJZ+rMm
NFCmWAnZpI1rIHGFcqGObrIhQTF8COSodBSj18pXSgkHTSWvJv2Xe29GU3BIVvYl82p3gEV50zpd
/yKVYKd2K1ujFpsAaaNO3WFhcWg0F4w2btJXHtXNrDcgTxbi1dXfeW3kS8InlvBndVXhOTxa8idh
xsEBBrYVI2GUkcrnXYWGOgj385dHh0DwRv98m6qo+yJnzIWDR4m2J3csm4u16BnfbUS+OchVDHD4
wseIfm89XBPG70RsDLtmxl6S8MS7tXzsse5r8l1cigqqoNR85/4GgWS1MHHVyW7xsZIS3gh9v50v
BQ0zW38xX5/B2rzCutIuCdpG6wyoC3lPh98aBzRRHJRbaLCtt9kfrWn9SnS58mJuc3iA/cRQlIe2
aKUpOk6jXziTzzU9LgfXLtGF/dHil/L0njAqEV87iCp4fd9xhvneqe+A253D1U95huozP/WbiE9o
BCEASU2/GdoMTrV2VQqBBJI3OIGIOOIt0idsqaa0sA2NHRDN3CLI1qSlH0geiE9qDcFyxIz3o34j
Hf24EPjBPpB2ASFp8z5q+9S61nKBuC+8fHcMAYFa/5vYTLAcr730HW+IUZnct2x0OBcbLLsSr7Nx
QAXMwHDs3dToMYeK9dhSa5PZTgMh60x+jvf25ydsTnni1r+xMp5FSQMYvNCt6GBKumiNVGcHsM6v
vjwUkNQgTfd2HdwbyGrV3otd4fmn6fXT9lOabx9egHyt10a3Lnzb4mQCELvzuQnyQPUYI1kbqIEH
GyQH+tFTgZNc63D+0sbIQJk9XSw42Wvhe1gP+yqI5eM3afWsM/dfoEzmY1vGXIfMT5fZR4HTq7pK
BG6MnEDPPeMZI3bg9T6y/3LMGcDzO+YBftvrxJ4xO53OjbtR3Hidyzx3tQfnVIJ+IYb5xT/IzfTM
V3sRnHJvV/6olC+URcs1q8YFEgWbelNmojxuDWLNeHDUKz3vbJBCxWpsJuDmgEzjf7Om6SmMjcEm
bgTWvgHb+vNEQSw3olWaX3UG9uPTt7mV6tPH9Em5eYhI3sP8FoO+S+WbRab+8ktJlUXCuLofDO05
LhnwBIY4HNujb55XtK50bmVOauypJgZbFBqR32tv/csggEaKsteXGotk0IZOALJ8NRMN/4R231nZ
SjqBF94xVe+aImMPhQlpnW4QbU+yptDCyDogJ6UbNSuJ4u0/6UWA6wBL5G0i/VXStzCxaMDaCUw8
s+e3RE/9u24SMQAOeTmG29GXUgla7MkJLPi337jtVIJJ+dhsH31uM2eul75JealupgEP1Kkl2E+Z
AHUaVQUk0zbr2VvKc0N/4djHKhSpLxN6QC2IBajY3phn8xRXI/aI/BgmkjxWCYg0kLBpkC4hbVN1
ELE1wGbBEMpLM/6iO4+PKbLQRUBgCi+1mfuNuy1N77BdYDurIuiShRxWn+Evve6ujxHOCZ7kPxCs
qqweSamhEjKkxzj+9F//IZgDT0A5KDTH3NHWWXdkSij/yYxfgAEhZjtiLDOa11jMsv8b+aUjn98x
QC8FjtE6j0URMy9UU1UhtkivZPcnM8gO+zxzIeNM2obWhOUmClmQagY4DeF2PXQa5/8IFTOAudY5
JE/ZIg8kekgXGcizK62TnMq+alMVq0a6l4ggH/8GW5yP0yaYPZxfl44It/prgul+W85CLzpH8ctG
/Y3fCHwoIEqusHA+9koaEekl/7sddeHHddJUhfpOmx4WqNc7M3xkWOdfk0XOdlttKxzUgXUwKFS0
Y+mQumVr+xl5l/sxvNLUEvR9z503MckbbxWEIXmb82DWjRZriYmecAJPitUNlSQvmcY4wT1d8u95
fItn+B7FEgqOIFAVATSnqCF0/Ozb+WJ87yPFW2QcMaF9kNPh1tF4uUHRLgWFMwsLsYR+uJkUzOP1
r/VN44UgnaSNTgMSvr/PccOwKwedR9fc3E9RsDvRzjfKPIzZYPUROXbuBzBVrR13CypIgxhLxrZ/
MFdCVgzMqvCLryePwBKcf1fB+tPOGITTLOvIDkghFdpJntCme3HNoc5TN9m0691XmcDcufl3Rzye
BXDZOnglsRXttnvbsi3aZyx8NBv6pv6Em+wuw8iA/GMClWGoT68g2+4oybFVxdrRWtcSUkC2f3Tb
9OetAcCDkN0UORKMs5bKJi0puWmQOG5URBDtMpl7T1OeKhysyTlRWABGFCxKtsOaiwqaK+IrC2hC
6kLmJZpCDn2hmgY+WuoWhnBsk4li0MBYi0F/8AT7OFquX9OaCUfHyhbRrgvYPCXZ/90+I0lYwm2J
fwV7I5m2iKWW/B/sDDL7ZMaIlX3HHFy8ckMJx5rlja4qe2rQC+l5jHM1GGNWHk52IJt3sF1IPWaK
rD+t7WZkJwNtpg6srs5bVZ+JPDZ/DUjGOVobI0LOAbAgJJJGwGFcpZ0ouKb6Fzhb4dT5E79xmOVs
37aP15voENg1dM+ip7FFg1j//RvVbzc64F+8g+zbgc4kcvkAqnjMmEQlIu+RN3V4HADGt+Q+Fljh
Ys2/u1pDbJw85LgsKqx7iCIPli7mJqeuk2ir0td0MFLT+nqhffzwpoPcoSQQLCEOTdNjfyoU5OKh
7DKHXuMmGEGcGpV3bdv2xciIGrd7i77/GKXQlY3Kx3pz9CDC/9AtRXrjJiwrM/c5IdkFRNpp7Zar
kAfvNzIwglcjoVvWYXK7bzdysEcyWRZUPrlfrWSOtmOMyinyk68hyafVxZ7fCrPitgMgbmDwTE4a
aiu9ozg5sQS0sa2ceIxhNB8ONOxsHbYXmWoMzevhte/Wyqhdz3sPjj8u+3mjR+an7ZCBylVlHHIw
zs6IHlauTwZw1PtTCraUCg/dqMkhvr2WStat8F/gto+v28GAA4xksNW0eA8yEmid+Ib6Yu2VN62P
qx0IuZfVdU3gFxXDKg5b9uPsSbSjp+lGqrv/YJNpp4lBzkuXwf5+AQSKhamNX7u9txoiaTOC3ZtA
TQzFA0ir12SN+DwseehvoRyVhYcHMm91Tz4JOZJGyJWEROD1gYiJiJDD4jn3u1K8ZvfiGPaxfuPw
huwwDhSRVnstJbAjhETdXhIYST0JmmwpMQnHF2aAWyeLm2bcfKM3xEHa+1ySq6XAyTWaEHgsP3bQ
IVbpY7xtpxcC3y2DNELEBvRR8NK75Bv89REsUCrpSks15W5KlfZ1zha4QWsSK1nTCvGtJENBqS/1
xWtadDXDMyNXh6vpl39GkQXaDXD4kWzmzHyBIeWfKVR29gutWtNVgkqjEPxgYRcCpz2l5z3teXCy
Wt4fSt+vueSEbQZqrA+o0dlZsQ9fjgCsVF9o6jyxS2w1DKAIOOICkMyYpb1aIqGjZBM07SgL4YCC
sncZOzT+ujr2TQNMvZlAeYPw14vc7a2/qkxE+601AKOgPtth+Xlozw5KXQatS5MqMP1Y24tIJ23X
/SnEtDzTVkEqGRPJ/VCD8mtZ6sLFsQ6Sjjjn0xIhWK3ewrDiPbX/W+uHoAVgAaktvUajQHPRMBTf
8hQ6nHeWVPpkEnclYtjlgiQ97Qnl3gNtjjDoLg2CkzLSQHawAXPi9i4CCC410JYak1wFW6dO5JQA
qZwOx+VS9Io/i3v2/VjNo49T8m5R6Jd49qpr1pxg5Q0mUXzeAEpBxzRGJBq9pXLjvJORzYeq4Gjs
Mv9d4hosNecjY8OVWL7e/A+QWIxBj64qYoJgZJoHqyFLL5CpdIPviBmEdOZZ7BT57c3Qkahis/Kx
wuO8Z8YfkazrAl2VpQ1AUjFuIPK14zzC6VElo2zWbNq+nTTqAXxftkngYzPM0bu/00PJ3fqQIGph
QOdnuCIH1omePtGbAiLIvRd3WMOIQp56NcBzPKOePnJ9HDTu/8svhCO/sXAblmf8CjnmmYibrNkG
/6oUGwUYjE/arkoEQfipDP7hVViLB4L4VbhJ1/VjQbDlfdkSBn79pcoCIlZAS5dOaUopXO5+6D/3
xsSClPdSdyh/vOUHCXMf1mmo9lYUavn6RH7lom7Wb3peNHrE8ctHcmzF6yApgxbwRcJkBoFuldqY
KOFBZ0zjtxcUvKZQdM/fip1xJkU04G0YbOel9recUQ4oYPT16gs8bFTi4fDKhdfSS347/958tzWG
MpnIiQscfuGNH6BrD3DGM9xrUAXKzckYf8/OmSci2xEHbSaOARbB4vnnOLYLdG/jQLtnBnsatVD3
wVip4Bv/n5q8bQ64vW162Rv1eYMazYNsrw86sVX8VY9xsq+D8F9bzMyc1ljZfape+L06e+6PBNpJ
a8mGXlYajnQJTuD1J2sbOK0L8RYIWCur8q1I+izhLGWNmGQtKai8PgxNeFfb3r64fbcgBsyXoVFZ
DdcAwi4OkXf6fbrRKAPK6r+Afek7VNi9IP+W3uQAKMpfpwHoDVZIgHieAA4c59hxOVUYfVXFAV4j
IXqaLxwmV7V4aNpT6dk6U3LpkiOF+hHx4nKIuDRmCQmZicHxYtz+gX++/6dOLYVS6y5Tepdsg7fG
8EuS2c6MMcMb8iPBA7lbcey0ny3Q0/Q2+9nerRHrZOJ4O5m3yoAitKQaXSLVG4CosKeA9LGpApaN
0RWfW/XGBuFufZ1xThFvGMCzAxTMKbksA2lGIqKLfTe65DjKEfeiSo7G4pkfyGjpeGYcsKjEDoYQ
Csz1T1WbOvG651a67A0jZHkMgrh+ZZEOg0M7W/QTq7qO/NFtq7Sk9yLlZ9tG63ZjRvbT82djALT6
fIzdMOV5yvsUNbURA5TMf7V4mq8REnsdBaQTB6Ep91ni/v4KWIaII+wDkEwhfz5SC1I1cX3E28DG
8W/yLHHjj3wsFmA3bii6wuFm2sQB1ZTS+4cLRcrIsuhCaA1qwuffym2qolCZ8GudSkOYxrFidfA6
JHAomMv2g+J/67eDM6N7IA/OduqZvJ27eZLdkcgk234HXSR3uttnniaN3k5qBVso+1aET+p/yFq/
dMJu4LhNg+fumMofz5e0XJMAbjKCqaafWFe9yatvUwgChkGjO+7YIYD841rcoQ+ZTVgy1hJ9Erf+
JR0/4FqEEuPdzFN3JYhbkiur0kDxq8jz7PKOYONZJLadHZ81UBurgZzrp3TSOuzHJe6pcIrMkFQQ
6ZGT6q7IgNm/Z/hMoF1uul4Yoxc85kA0AKu1tXgvKWZDQorhAX2jCrhsxvkaYXl2/bbRRCW0CZwM
+csb5SbY/dnU++LuSGvKDwwq9hOLWe7qn/Q/I+3aW1MbqfD+E1DVcYOkoY4UY2u7rui1q2rp4AQb
wjUbh+rCZi9EltclGPRDT+XCIHf7l8TTkX9huqCCi6l/tGjrt5ft+lK3TehUn313tkmsFWgoYb0X
ChucUyb1mRbhc+lGFAWBrg4afsck5oCFgRx0Y3ca58qUJMDfcTjVoipc7c1MF9e6IfTw2Cn7jzlH
HjD9bsHHvTucrJewUM1hJ0ggGG57sHJt+AnkznwF+gmq9ocVqHOEf6ukgT4mviyp8tsfEeGtZCxv
cIeGxE3mE0Y+YTNjjezSQ8/eXo4GyDOk6FQULB1XEO0J7F0K9V8suhkHxLW/zaH6KuWGBKU5tGLd
9uuUAQq0g81/ym//Qyy929DtA18Y18/sZhPaXeXdmWMgXLuVO8eqnQiAjB2KWYzQgZJdiy+yy6BZ
6GoLPricDK1XQ/zq1Z4xJBlxfytFPNN6x7SShWhWfGq3vX9N2+xE0l4WWPsdA/Hzs3F/O5voo5h9
yMcim5M7hhcHY9N+uQovQt9RvXR6pbS6aUro+nXhyWBRj3k4zsWoHhjLYqSln5oRtw1yTI6xCgC9
a+kKV4hP+nI4ND59MEhhdzzDnW77YYe/YMJXH5KL7k3YqpKv7YF3/p8/h+9ZSPAnxCAmmfcrqsMC
GSk7aINZV3XfIeJGeWVtOrod9Uv/6tLS1uBVu2D5GRvU8KWUNtH82Bqg6udV2LXyVGY18tGj6znw
3+uekIMS3pD9hyip80YQxF+KUFmS0+Rv/WCFZR3qXRFEp0HeVgWbpujRgMap/mthuGjNRnSYvZ8F
1m+G834xlieV2VyHs+HN/M/4dRiNImhw0dcF9FSIhDuVXI7AGka399W0DGDGV2qL+FkB0u6v9/9D
pGqBolgZwz+Vsj/O2y6BE8LXQVqE7kJ1zANy8CIBcfjMPnm4f+8Qm96lK3cEY0Hs3+uI2JxogSFj
UbHfVTDPxjobgOIpkx5uEXdgjSmgiffO5CAElK/ywShN+F95lK2YcBqzMnKK02Wtb5RK6nVG9qGm
/cKsF/tGbRsXRaSNyVoFwG0JdE8a9K0pfQsgTeRuOUcjxCkK1RTljbJRqXEWhBdjmMAash1UCd9S
KXQv3DtgtWZctVdkiDUDE/lorReyKjuyImn0/yO/wqHH4HjIKAG2NorwyWPsG/qmZItxmoUZXwdh
QH8BnGTZ7bxO/XeaOS5EO8uxBuVKcykwJ+cMqNOGJ2DH04FVE75J95sn1LZDXEPr0fFK3vNQjvoY
qnGm+lC7pRoNb5x92QXrizqO1jz2SqRzaxzW3sqwvrMUyELL91c0mf66aV6kHK5ncmTyd1Kd6apD
EVhjx/ZLzfMuGCnpE19Sw2cxpTTkqyYs9vc36yxhMT9SzRTB6MkL6XY9ixobZHfPd0LiEvpzqABM
vOD40tBtPaxlclpX3EBfG1R2ev/ePW9en+dCHTkJ7tjt8VwwzfKMJ4fAwzLFIGYcbLfHlV0sXFTB
D+ukra0M8ax/KrQOgDiAhqNky4ztxbCUiThDX4bXObV+7yaYW741qE7hJMotS4BuUVgcGRZzPnAu
as0fv1WPK4jsvlehnR3GFryy46nd9g5VuQBqVq08T3Lf6XPunmqwYOXnV6zrHYmG35JqvXyOaiKT
K182WRi/VAs4rBGY3jE2oPmbEvLwS5EdlSeIBmhPzdk1hl4dMpD7Z0X7zxrSaBu1gVFajCT9U++G
KBbR2ZFvTVVKyQ2fvbiGJe+PNM+zfXbfVoM5WDxxoWRgkV9g9XHfNfaWA2m1fU7h30Y//oW423ml
z55ysUsau6gG4zH8xLV9iXvMu+YrvgQQlbq9UF9cFgZptwkDmc8rSMM8YJlvtOx98fecOyQ4Hakk
jIr4cMrAHJSgNfIi9N66GO3c39jx3eJH2NJpZXv8rthYfiWlfQHam9i/Ijz3FnHuEAqbxlt69Ohf
rbQbweGFo+i+Vm5jkNDLDPQZ4TexbQtsrVMoEyPfVNynHwRhpT4lhnoMbSmfIChFjOIrr9B8NAIB
bf7XYGp/WB+htIA7M792cHTcExSR0nvZaFF2ayoKQ/1VovSosyWTKBJVYtfbQrQ5WNXUAGFFSZSC
jruDYkr+B6Xu7j8SQ2/4bo7xW7Ds5zVq+e56YdvZaXJdqgivOa0OVk3AVmbnrcrn4xXTfbu4DBJZ
o6eYaj7xZOgSTpBi98J30uzIdcg6o6bpqyqSjBBK8uNFljUWHqAUq5ydI1gv+w6VLCzz4zPp5aB6
q6f9v9utr0lr7mHANrFMTnOqLAbJpfbABsjGch/gsgKnlKI3HQLlNLi+KoqutgrqhWW7O2LWsTtT
jvxo2AKk4d1B94e+1zA7qXE/R7tv1BpSG+v2j4Ly+BG8E18peXYQYYqv5aTrw5moI98lXQZOq/h0
zRGb0QLbtCoYL+7Bq71rAIc0RHkNowN9eN1zPAVTUiM0E50WYICRIwOMgjcbwTBVNYtfQEN2QhDp
gERprrpBFBHL4Z8SCDW9xL7vP8cpLkPtrfOI4CfPmvGELgwkYD53HLAKHUWMZB/PSBGi/WJR8Suo
b79N4d9G+xFaWszGs4PimdHC/FomhoFFf0T4rObLtkDQKJaWyeYJOP18+wPp9l0E+kflksfnr7Fd
YZoClpTsQCyoq8J0CxUsvqM3K1uzLE7XjHO5pHjaGTaq+EBRklsvlKoCHCz8/a6RtesdzZ8ridQs
HRY95N9Q07dIAeD3QQTmVqk15u1KybwPjZu/4uRYHItW4i/zgGi+TMyw9IPZyNZwqWOCiCAzuRlc
L5X3Xmc93AmCkMYVqNRLxLRxEAGmDdPdOkaPxYOVwxHDG/P9vDsG3UyRsJSI0u29dRFqgSonIrKe
ttRmPI+C++26s9v0zCaLRGqOuXUa9EjXN9lPPo5eJSPeuOKtlLbnfGnpDqINBFpXBtG3092ZMybS
XEC0BRJ1vhaQe1Dt5axnIzpCALV5sBT2nmfjqaYp4XnvORorE5D1jqUqd/CWPFJdHIrOgwith9nB
12rHbWGBeVGNrVONEbO9ObGW5tc+eTwt+0PiyBqzbGtuVMQx8qWXxlMYWaYHs2MoJucSD5MSyPnE
BW4NDdts8GFQZvYcDk8C3XkUg0A5ccVV2BXVVKCX2G/1Z5pY4fS9s8MMS/LSoOI3GhGuaObnPOhP
ebuehdbMH02db2ju3r/dYjtsFw49WorEOeU0r9+G+Saf4iayAdWZIjZ8zdUBIoYv9w5rzBcJfGXP
V6ci45Z19xOPgleAvZgtupazwwRQ4CfzhPl4Xzl5YHGYZelTSyhbJlleOePDLuHmDZDWtwk1Xiop
Ns6cHXZgzZiTdzy8DjNjl6zP1nHFffoa5Zb1zFs2srrO5kFagEWSorl4NHZ1sl/CjELC1s7pvaFY
ERmkrkjzRgukpwrDn45WgJm5QSXC4Jr6ppQsX96bmwjq6rlJVvACVpCJpRLC/MxCu0FqPLHFAeMG
FSDXQrbF6GTzi5ggrnB37tE0Br9Qq9KPLe/kQHEapgMsuOM3oKd+esVHsTiwlzBCjUhBMiScjnaa
yZ8IeykzX3dcgf0Y1cRgqxZp75m/aiZtW2rnDQBvI1WU5U7Rm9/IBxmmk8H8o51XNYk8/QRTDrQ0
3YWIBQEHuJ+L7SVKo/NwsvwWkm/e6w1M/W3qwL5TXBi+EqwTpW8v2IMCEf5eD1ZOifhfD387DWPZ
8NofFpLzmb6G7PjIXMeF6sd7SDdPd5jLXdIPY62VLxSngWHwt3lrnaA7yCnNpLb5nO0L+PStDclL
e0cXgfSTtuLaq5Ab05+lHS8IMRgBjsUXU+qH0kc/++1pU4dcLTIpZkhCoLylTaHBVKQxFSkW+hmv
eFh89dpTJ/0Q8XFhsJKGOOT9fUwxieJQctY4+a3lglXsHeSjoFbmNmMY7fwl0abXdNS3upy8J4T5
Vsn8XWlGfK8tp2RBrvMXAdT+yau8J4F2cK1CJ8XFaqv2h7GankBEpIGIXYb56pazDrwPBe6MiVwy
AJjqwRz+xc4PBzfw51yRW1btOWSHgO9DFKlX8nwZ4Hw/KhIjoDZSut381zsdp9qq6O8CBaHBv4l+
+JA6Gav26vHFo4ivMccxtmhRwsuuk/1ZS3qckYZgkUgqSLpFGTaepeQRsC1PfXlCJJNnfIU5OsuV
hR3Cl6RqzOrj5gYYkwsRwSQ8ytIAr7lQIZ0pkKSiPRt0E4LLvPuYijvFFsxZ/usmzYEpFDWACPpD
7iSNUGuYk14Er/kFiExeyEFdNyCeJkazm76wcnlyLGlxM358GMlojruKQR38mwo2dVDKhNmakBug
6bGUgFx+zTWaKyxhbbeHeUjBfvS3YWHzwpFZhJMEepOzXYK98mw27YV+kgs3ZMQnNYPWpmo50u5U
hMuP3uT6Oe4rD5OG8RVWbtUL36mWgCxjV4QvWe/qlWyXH9mCMT1IgFboJ41561/6fJBjylp2T5mD
+LJ/875tzUxMPFZrhMGV9uMayFSaWnZTa2Cng7+8F4PWRuNjhur+JwYWOA4Bm9xL6EaLrYa7ZHwb
RFpHATgWK5Funr5Rc/JCHz4i74uiavr+GpO7h8255chih3K+0fEDwoJJP8TMxPJda3Rf9x+2WJx9
ZKtS0tt/9bWhvft6iMTjhh177aGyc6zxse3nOwcS99Pnu5XGV/CJXaxTqId5FeMhBFl7h1z1gM8m
Bj/SZRI5662/zZ7bgTJ+7IcnxMYWJZnjlNAeY/2Vlxv0wJ7Bcy8zf+99yi+DEqPwf/nJjaZp0frm
/HtIJcvjc5C9TIRkT7zIP71Oe4SusAhhlYFr7Q6BacMuRjOybUO/WNeYGXAnrd2To2derlN09TM9
fUgKOLLjzWsr4bP3h5Ry5a0wXgVzZykwkLWqV0ZBhdt+EsPx6hUhxApPmwQIgEW0w7PWmfNItg+8
KklKgoDRDqYnzRVfQaH1U1ehHAfR/CiZK2gUxL7p7BousW0jQpTZi32mBiHki4wUrW4UFds/+AT0
XPS0dC/2WwyODfbBBw4YMfqSyMdQFGKKxK5W9LJGrjUmlcSfpUqPX78nXO9EZMcqqg01uL0do02j
xps5dW6Tyu0VClPj6CmUcRCyMoVuQeiRsUcu/t78RM39heVyLsrn6+GlgDOV6lzo8In5sRTGibdh
ctarGjbA3eHjxiaVyxaqnAEo3JQwPeHxJ50rsVLul41EYSc3bmwEMdUaVSXWXEzz90XLzrPsVq7t
9qFNxhtAXNbQZvYhIrBMX6M3zSKK0cTKgYu2+H4+o9TM94h5LX44w84i9eqSxkzUHcOfRuw4WZ3r
W5OorzGGgM4z3409yA8OkAI+0RW954IZnRZLG1Ct9qiClqDvXIm49fyL7EM25nxiNBNEXX/Xdcwy
UEz1YRXokiGCiv6EqdGES+7xTfpZHAMVwkbpazJ2A3fBTxg5kjtCrwSyZuWuTo9E4V2SaCdHEW/n
Ul3kn0S10YLBZ8OpaXzBs+hpMMSrY3rXcld+kr8FiB1wNQyjoIcDl/Mcm9+WIN/5nRkBuU489LDO
GOg4GFyflJRlETnykV+JaGvxXFGh+A+zO0uqia/qXSgjk1YivFK2rEef/m8C82wlIE6zF7Z/mojN
EOG0jw1y9WQ0i3v4VOk59B8z+ZKDUjw8cEHN8TPqulPvT/ofFlS3RXgjHIrxkkImEZuMde93wzJy
HoMqkpbgvMA5ZknQvjvxzitfRxJ37sP6UXhvFyfFilwrvMTwbLXiYikdWU25uAjH1j6G7gswIFCM
nCrjxFGG/B1hzReF6Ftvymnotlz8CKuelvhpqzJ1UxqRpPQ/0AOIVJ5IZxzVHuB8maItA3hKWZ9n
1E6cDF+gN3CVKafigIS2iAvWsbzyasqoaiPk4u6whgt7gydLx7xWMgVuLtxE/Tk4H8gbXVbfkSbM
8XFX3XzzhB8OipHWaPWgNrE5IvjLzfVvjD6sQTeV3qwps+aY4+QGBsjgWNiONjGdMjqqXvWcvlcq
l3OYn99pwihz5bVXfl4JQDmJFlzv15qKwEtiD6IrgwK4S/KWAQpIpTCUSD7tx3BLpqqu81an7JuP
iVFxgDUaKoy0+cKmiavMoDVaFg2UQZfQ2raWAWSRJhxrtVC4IVGZ6iOPaevaYm4SvbLaEIL9vwwV
OIDXa1p1Ipg7Sf3VjBWLI8cABf/CRdsoH6mhgRZMMZXzOdQejI7RR9gDOab/AmHWjU52gRfrCI1S
G8Qkn/yjftw2I0XfwU5hzWqzn+DjvosAM2QMLn4djWPXwlQ2C3WJqYt4ULag8L2oEb5gNxRQPmdi
DW/yzTIy6DLJ5qzWatXT1O5JGsD2kCOIEUwAfHwUr9fOtsDN1PkgvobyI5JH5BBG6IVZAk15BE7D
5PGRmK7PnQ/yy9RAweIi9kZ2BZyyZYii0y+dYk2t77l3JVIxkDWLigq0c5dbjNeK8QRuVq6fGEtr
W4priyF02glmTpMQvyQLPb2US+tehI2vsk3TUF9gL7gHKTaL1TlUrN4kTdp48xa0BOdhTJHLAAww
XgISf5FCQkOcrhT/7joNlrtc0tW361hoE3Loc5Ma6shTtRkz3zgCx15QOdJ3co6I0sQ5lVR6kcQ4
yrBo3H0pLQDrMRLoSXKBP4j1F1Y9t03ozoq4RZsO+/IsYU8+kNVEXK18B3iKSlNbjMSmZe5pvlAV
BEqnRApsEyDRapKYdMwaTDEZ2zIoUpnWluOx7KH73pZms4Vxow0L1P8qWiDb5MaVV0uQ7MRUSsk/
2oXH+senZivMfiCuLVv613ulI6OdE3GK2Y1PsEFfK6UMSDaolqtuqqrNpRiy0QkNYdeNjpuNviUP
SLfMmUoEnMFk4OqQYSa9tQoF0lDvG8SE3umU+/tkl1634DAVEHYtJOeAibV/aTCu8/qGhv2hzPvO
DEkzL19WKuNf1lQ0ZnWKg/c0N9APmJ08NKYlZdgDH/z6QnAxdawmiKvQAc+CHfSZWs+Ht4xao7Pz
eyYNMiH9cQQ0YocoLUW5Pph+9wWXMv+2S3ORaaLf5IK06qQDcgPrGcboMTkcebXIBijSGhFPZ42x
QOw2PCsjZ5op1T+2Z8yAPeMRFqSe89k8pa9kEh+ylfvu3YUIMRi7pJOyRykF+4v4YHHqChsIbIt3
GqVxcG9p94jAZjq118zMLecoB1F9awYDUk8mraPKkWCWbhWgSvmDU71gWH21jZmUMX7s9rctde/8
Y9OtBG3iwGiSPNW/4cBFj2TSKniRzQZmEG8qtOiWzjur3Mzl/t6fZu7m7i8Sbn/bxg3UJigMGss6
+7sflt1+Lq8cBUFA5KfDdJ55TlhYZQT82wT+CaDPu6/4/Hg2LMZ+t+efd8TmCA2XmAx9x8vn3O1j
Oz+Zm16mG6Ky9cQlieXAPWd780zT25sKtoy7sy+UJ9yOcydZ2rfPrgux+CgpybqkqR09JVoLrtit
oSMgWvix+D9h+iI2fqYjAYT5/+RA7NnhJxHeWjnmP/lfT3w3oRRLn16uDra1UXHald/njtbtYUO+
WRVcFrrOGAwOe0AnYh8Wom8nOr6O3DtY6N5J3ZRaHt01mB4CjER/qIV2yPV4TeEO7ZeA85suOipb
Q8yAb5kXzJvz598c71GVOf06knhZZ35tqFClxCD+yuKDeBa+fYiNFYi/WAPsd3Dmht1DbFEun0I1
VCDPtTsfJprfEXLrAkkT7zhvMSCPSntcPPWJmaPRprDR9Rp/E8wtD8rrDPZtrtoZyK6KzTctS9PP
PkisAf92zb3AystjJv5w6Y6sX8xG2grMisyIfbIxNYn5A/qxuS5FWefQAVVTM799Ts6Mp98CAFcG
1WqQvIdR3XaDH4s+LytRF2uERzLpd/ZTIC4AAv9RqvMbsEeDv08wJjNZHfS326kdpeXlu8KYbrDb
IBe4Mx2c5UA/bYil9CHindIGZZJERVklopqZuWan0IFQ5IvVBr+EiW/OkeHccnQbu4DCvUBUv16o
aaKXh7BMvxW+5Sa+GT3rGVWYWM8GLqWlcvN9hwZwzWXjPUbYV/O2OD7zPsH4FlxGTCGOLqrD9quW
qJFhLHYhAyCyejdZZyelSL6GAX5xRcbee3ToTUZPrwCMLQGIbHFTsRixVd6EaTGSXip0j1nQN+tA
5EVOmXWQZwd8RUE4SKPFiNEFCUX2bPqFhmNDeaLFkHt+gJfkq2ZxWQiytSF/Rmd+y1QaSTCQ23LV
ZjqlP1PC03LW2jlFAsfgv2sIEMX8gWf9Z1u3KEm8J2aDcwJmmnp4rS7Li6QwcldQJGTV1Kn+l0iV
yMKBlmkMH1hnC21lgOghBX2xO5oqGmMOIILhh20GUY0FXzvR9VfuXtX3WTKw746Y7TrGJc9ym5BL
R1kFFRXYB2T+1HtFTIPdtoTmf/2yWy5+0jc0tsxEz/SoyQFx5YTkQUYyZY3nJnLNLT3sylfIAi5i
zzfP9TcdN9zS96RNqFtPltNCLLW9PE4kB3JH+aZnHI0QKXsV9SdoZmG/faPMkeGfTXsaKgvQMOI8
Btx+erGKAxmEUSooEfxFerkV6ZAo+jJU5R9yo++APS2FMcijxWbq9tGEB+g0Ig88ZjQOvQ5qqUbp
matcM1o5PPHSFnicYma7I4/BhXyiRyzyRR+XyQURmrlwZ4JKnjZIyINJrl0O+68If9EoMVUvAPg+
NPecE/kX69x/+FGGU6Z0R/eDZhYm0xJvPHhTJQojWkzYEaoQxbrrT0KMNkpaEaGpfObTuCboeH37
0ZD/aTjpHhvkZPF686RA/+EGBI5mzF4fHpfSDmQZdlOD0LlB3Dww2Ki8bA1B9UteJrQPlVpxRsN4
03n1MdSWG72O3+YV+VjAEcyIU/08/7F0WnZQYAU62jtB1SURj7xVKpuQebKgvgzkfLQvtwg07tkS
Pv7/XuSn0uewmxeR6b4mBY7d6yyt215mnhZfr6zEQgTQ5cR89XMBuceXnFMyD31Khi5703VNhs2s
35im4FhYYVFoSrzssfYbDgD9AO3kpHU2lawZjod00clJgxAfln9vOcStaQIUutSqFCHXbkLX1psJ
eVcXVHExr0r6xNEHuCmK3jLlIe5oStIr0M/Saz2GFPjAmc7eSUhoNllmTzKv0slVfUPpq+v+cjWE
T0+1vuHEoUIEkNqQEMui4qyDOB0oGhyXptz/Eey03jdlo7Tlwn5QZWKQAbWVVZAZBrNiOUh9QLU4
qysdNpgrFu2ALkYcOhDueO8wz4ntUrWODITb3hJLH1bI7QB0COBqaKrPXVB1ItS/ecFXJXJ28im+
wc3l0zwZR3T11UlppIMvvN6xb5wQEigSfVox1B1fIzOkzZoLVZ/3NR0swvY9qdxpNCgFYhZtXZOP
jCO46BRPSKou4ToJ52HnJmD2RpXM0uu+/a5zEkfakjXGqHTtRfskKsLPw5MLBtTD/E0AP0UL1zsj
AnCCUW3ciIB7D0WqR4xafTwm8K8tpEvfRSWY4cP+eq2yUSDTilQxrR6biE8/y0vI0kwTSKpy5Ll/
vpVMvtDVAE+ybN5Lfm7aLIjgCKGDtgsW0z2lP2O55bV9EmDMc+RoaSaaUEmDSQ72jMh2LSt/B0+Y
iqPxGRbajUqgLaUYsxBy4cOxjo3G3N3CkBKfZWg30+9EUqHNPgu6Oek3B12D6nQxkWGzEGUIsWWS
aa00q2UoPpRWIGD6PurhUSkpeu3KLR1dEg40lVnFpjaxSwb5WctUwWkyiRQyNYX0bWIx5ialpc37
aQdi1z5kJT88gLdV4vZlDVl/AijYqaebmV+1cQBw7cuc35hFIVgYLthRWqB8/C3E7n+KoI+Zy8CZ
vbFXhACSsQZONBTZusePXEl/UaG9ZNY0bhawksz8sQW4YNCP4QCrtN508CchA353fik4FblGN6md
JOkW5rZ4hOzfVsZfIICczr5pzV1LYUT0WsF7p3+8Ojpu3p1xJdKYsGqVWTY1jc5AULkvMjL9aubx
H9A7zTxaPpKW+2vuJxU8ALRhbNEHP3THiJG0GbYbBv/3cpg7Sa4UfxRfx41sMdhFY7lAAAWafpn/
xxCAbZkD4nNwIX4nQjMNMSycRzHwy3Cp8YUGHxoAJoQVedDcnaAQpVqaWMJnAxiyGctBNjDALgyu
OxLRQCl9x+y+WYHmdVJK06NSsoDMJb2LID5OtyKIpB9NnZcT0aS9FQ2H+MfLb0YkX4ffNo5bYaSu
3xyOgfCpBNeId7ncK2uiEXErT49RliIaMS3AHSidW+qcV3a/IFtT/6dqQkpuE5qCuazeQswK6kNM
hKsP/x2gbkxOlVuZwqbzF+cJtbozllcvX3UnrQDsjFnlpyC6BbMOUWbJD9GU9/E/DHqkQ3MRFT6l
IJMIJcGdC0Ec7tSBnAKroVR+pF+hPtwMowrg4nQmaGiCUu+jT5Q/tWu0eX2+az9wPdhQhuPDdMeX
tAwud4tzTfhmCPlcl9aexAm2GPS2hC6OnsZ3mhTO3hstVrKeDbdUScK9kCh/BM3EAlhRHumUZFML
AQZHc4ejVP1u9RyeI1FNmt3XJKDrWFP40TxaniQZ25Eo3ne5BSE6F8PABYPxKyd9OBVijXUGAKAO
cYlO5smVcplnTyZI9Xz2w4m6LU+xW8Iz4YunhZQ/LyO6ht7HQmGyfbu03mhkRrbXoLc/0DkaN5Y2
f88n9APV6MZRofx8ocNH/6L5gZIgUdGGDsvxQG6ieKToL0c/0E6yHeOmVR6smdR/S9XAple1B1qn
If323h2l8b1jwo4eegDsWKg/UJVpIgi4MmJe1AC0Vt/YgHUQdWW+CROMTeKiMGm+6YyKl/VnpO24
Q98u6B1MQyOeZwUvwbHobH/XYTWY+xE/HFcGOn9bW9Gq8iwDOwFWLjiXcCoJ4wJJ00WTbpHfDNm8
YxUoTrI1IlNLxc9lEHF4g+GiE4nbqoc3ptb5znTGka+5QUjbTwc7AitNchJmNJXrSICaP7qWyT6a
JfsqfSJItulDo8TtJ5gDjLeFcbl0+ibulJ/+4jO5u3ffbg3MnMV5SH8EInK/Jly0qjk0rsCCtGKy
Mt69Gknhj/kx1CInH/ZFw7klUnflbJH7mE0Fur7KK6mYQCIANE33AAUBTB9MUPzBxn+WWl6N4q7s
5NT4gcwUxmlaJiBA7CJZBTkyMLNEX8ST1VHXrPjSe38oB0+SNl8itwd+PryDAkSdbaciVIN2Vl2a
VqIFG47WDI45U06wgXG/bbNh3g7t+ga45o3BWALEf3572mOmOYW8PS2kOfoOH3DkE/TebALFsAAY
FPK3YK22OGFPvlUTMYMMlez9fzfV8LHcGnyLkIxiVxzwVAWeDSql6nv7dVAraXSgRV2R1tuQZFwu
xxGuO77f4k3uLk4v9MbiZyNLNnz0Dx3geJSIJXRWxJNVJQfdHz6OHzqeVMafhaK/nx3+OtXIbkHx
tzQw1zZvRo0UvD6uqC9VQOdQDtsRE3gXmlb4loRyoCt89jYDAUbSrxOP0WbmLMtNSx5PJlLOin1d
4dh9l4atKSSNtaN0ac+mGXNTMnRBnVs+r6QAlneG8ZnfW1pz+jwKW8nON9hBPnpi1Dn9ZKWMPI57
S8Pn8bb3CHDAtdBhIUIcPvIneoNkP5uh/mYsgvE/F46FWQWB2q9K5eu7eK/KzBRExJuOi18Jf1/T
mvYHutjD8lWPxJS/deEU5lXiCRTgMZ1kvR08fhl2K8U13mc0YwB0ReH0wOhJawmT2CoeXtWpTNdP
+6hICWjNi4XRCVWM6+S9VluZa9BHHEwpkK9TKG5jQrXizkX+pYu1ZW9x0g3pNHpkZFRv7ZhtsvTx
c//je7JDaZkFgZ+KccvkR+C1hqtFkSFdjYd8faB6D0dEByU3zVrWD1iW3+/cFTvjH1B3rCMlwoSF
65bGKebzwmI/HEOKejSOYxYlLd6bqAPw/zLDktx8CQDmiM2ZPcWyCHJBq2LVGIwRSW0QFG44J0XD
DYQhTZEwFG4vH36SlW/fsg8A/D+z9tU3c/77ufFONPKgYlkhNHrJEOyVnrSj+rcRkMdvE3MGlm/j
zJh1VWiVdGUrOP2L1GqIxBTCc9B101u4L/BZEyuZI8bnkWYGXT7NB6rM7SQl1hz2YAtHwZSkvoaA
5+XdZ3XN7p+Y/7Ojzt+Yv1SYBOuSe51M0v5jG06hIZOdZ0z3utKYeuRMbd7piv/7YnE7mFwJfpaW
L8k6MyEqnLy12HFx7rqMi1dIfY0ore01zK5Aums+5hQeh6pjFIK2anOnLNPunflvhN6aLrQG63re
O01qNE9bi6BsxGdQ8yuwBQpJGua91dO3spbm20ghV1xxQbmt3IpJ9dh5+46VpIbxYjZkssLU+6qQ
9RjKvxfVZ8f0TPP4nZKCDbenfYWdFH7ZAzT5bp6oeRmO+R5e6LYghI0k7cTcUhP2/yxsWFDFYO5M
rjkhBJW7hsTct5w4Re6+osr8sLNZtXkVcsPKUR/emyJszS62EJIF/V+NABojAxCVzXUUC1I2M+4f
NEarr4H7q9d0gK1vTb4MQJb2dz64z2MQX/w/DrW8qKICDOXj7yBIrjq5qRLCKLTSlnlAgtYMunzZ
Myy1lHjsF6rJ8rIrIa6eHu3VJ3ntyPCt60wT9DIL9QnIdH642C5HNMdr51u4G2nU+As719PZtm9h
kH607a/px297RSyHVd8mzDIDbTZJ7qx7rAU4FoyPPqk2CFiDzio+gi0n+QUCTRBGgnpOqntA/OPj
aJ8R77ssDHAObO66mdkRUS0xQAJ4nLmr3MP0JxH99Z9YB1SPtPhXosMUanYyJkiuXsg5+fzUT2vE
ae1g6MTjI9ZEO7FUYjfGqtN9tlvrWWi86OBxsVCIEzZ4FT/fVKX8yyUXkBl1kTvZ+K63UaHbO5hm
tHfJriEaZP3hpf4jCUQoCmDQysSAAz4wKu9GVA7baODAzApHuGjCZCZyiOj6SYaWJsnVzlKc1HYG
PnPlLOvlZdL9lqB7EudFDfSdR6dKt7CQjNLjGeXTUdsKaCLZeYz0VhbTtXlSd1r7vjez2bjYjDu0
fIgaJqhvFS046L8d/lW3mL09q2NplhQDVgagw2JdfO88P6lY3j5d/4R4wswvur1JsH8wn1fdrYul
GfEeDqIZ/BcUSltVOiTiKxiX6tRvAt6wVbOwnWZYUVTu7NGFpxDWA8YjBYkdAnE5taZQAlzCH3UT
siIc6+SzKaUaBC5ketIKf5C7u6D4kmDtVOB8ikisDLMW2VMG+oN8VY4zAmLZLzSmvqOOTcRfQsBQ
foQW2AMqEtb+VcpRGM49oPGBXkn+B7eKW7xqVoowTgrAdp6ZjHmSb+HBX+A2bV2MuJMeR1ic40Wc
eQJzC1q+7wNU/ha/bSvNQRafC30nhH7TkrmNmC62Uxk3mb/33kwIbotgUa7p8ioipJei1nrxt7m2
TTR3zkLlEV/jtDY/F71CbXnd15gbRz2K+3x+3k6nx0e2fi6+kTMJtZSiq+SSIX6vot6pZZYtSMta
yzILosOGEMe0NDEVyeegtQUKK5hrDyTsQxfNEbdV6nKkkfDHLfTW9fsfQ1yfNQXFfiMdfcD0+D7+
OgrowJy4Qmxm9oVv7lglkGWXrCUK/mQcP7Rc2WKnUEEUFo72wajZgdYA74C3eAiOPjAxV0M3msaH
ESrTl32TM5UCSgGy36DjmMAiq1RcJmnzKN0E7THNHGcByPWrnY+xuHeDn0bB97urKPhXA55V4eW3
CpEznTzas+P5AQv8KN4lTD+vzR6KCryv4wBsvIdwrv6m2SUaVz4ZHc6kPsYgUMi8BzVLcva92luN
y96XRO41dN446K1n8zPb8cFUfVMU0ZfhHepL0H6hFhVwljeUGYc0+RiaK1JwhymMlsKchsMnvbU+
NTFuaPs1n/AfUXv/WJ27eO1k/JDWG/nIn2VvkkIXtzW6b0G+bc/XI4+6T/5MJg82EeAFsTk733b5
ImjyOw8Ta2ouQMErVDxbz88tcGO95SOMjTIzGk7/oQPTLxVbh6XMrxNfiVtWPf4NW51NFL50xX+M
zKH4otQEZsqt1c9RiAei+77GM+vMfDT3maP+VRBnuJfD1ztkIv28+k2w1Jf0so3noWczZ7lEKpu4
0gd+mhJP4SoTY0U8I65V5HIBPHKr8VHFcaqpSRn75u0vmUZ7wibyyXOwpqX52Y8Yn2qNuOeKNl9V
rERQubHBCGjH+7d7xa8C3CoyqarVbiIvacqubIA9FXIUIZ2Dy/g0FSrf0nB6jUidujpk9BZwTGue
mE2S5dh6Rj6Nv4GThaaO0a+NYheEasYSeeQUwMZSkRgACcQHaL6Xb9lCP+SdarThyliHgaf2b9g/
EeFgTVcupJGNuUDBcqO1hU26hLt1RjqdyTcMCOIUKB8fcVRH6KcKHzKK+vSXWHCTmAYitrlwEk8s
zMdf/UdEGJvGkGxDnObSi6LxiaHh8O3qKab1FOVQnVR7GMMJWP+k/s/AnYZCspZseSN9qcBMvmhe
OzGBTfCdhNYixx1cHMwR8al4Hil3jeWpu8ZKA8Rsu9eTyPJQP4bsrnFEvCmscUDY+p6DW6z2Zpgz
qeH0cqYGAv8AAIYMAwLPWD+HQd9Qm2Sw4SYwKeygHAX35czi/VZlhHyJSJOCk3xNM1ieCTeEuhS8
enV91HI4GEHNQE9ibpuAQl5JtwWqrnpxGlCve+hTcIh+PM5hEo0OY5pLjuj7m2KiTSobf0KuCcAs
ATIv3fLL2q59bgySYoKo5MRbHBgtU7JqGlFC1tbKavcYu0qpIgm1Tffb6RKkXB0Gv7ZFQ0PMjdAt
ifWObjo32qQfBMTozr+JcgL+FVmvq1gMUJa4mV+afTfSPAAiS8CtKiI+5zedxWD/5j6k6TnzwzTs
nCg0xyG5+QQd37g4eyqyj2EihNjGjFp8QKJ/gTjMukbv1IHPx5lTJZ+5kvOfXp6BXXHPVFvf+4yE
G8BiHwAOY9BZZC8XdDr7lUKcNgpWtAEa598rfT6ETpSUBz8xbZMUjDAtPhzU5fPxCpxhUPrBcTO4
VF+c40BtSWu2N5hYAyEqZvdv04MSSZ1bYYcaeeFrK3r3aWH6iF5BtrwU+caHDFSyOEF9ijTRACAa
nMnjaHDrumwqLhq5PIBFBZiQ+XTnoB0lGLHm2YR16VRq8Jq9s18pKLzLhD3TCO7MBjFc7DxYszNi
RiK8Uk29cJHLAibsAXh8ly5Y0EBgeVQbvTLb1xopRQazT5ifqqig+eZzn9ZUi9Ue8Mqaf3fu+S1N
FON1YhaRrmt+nMKvciBuICl/vDdkvbgLbZ5FDH0tEGFpXxYezYLPryAiVkkfx928O4vsduqOwczo
Qtq378eBXIAPzP5+rUppMrHbnSP65/Rn7s+bbSVQKOH3uMuItGwhySb/q5WzGU0Ji/cQCjc4KtqL
gZ5mzXR01YUzrrumkUYoLj+iDLNTyTiQienyLeMRyqoZ5FLuqOBIhTdTC8CFOvRtY6Hk0FRK1KIr
iU6rJn0hpESJ7FZfrki3q7PMzG0rK0aQr3VEi7tfsqVRzac/ld51Pp1gOWccCRmgQWFLixsPLOCP
j0DTC8/XI3UcqZgzN/PlHLLWiB64T4cPPhcrek1KyLgJREQlIyurt09chBRs7WEXCDWwMdihA5sT
PCtXVMQy5iziB1UPTS2gsVMxyqq7ePJKIMAqdFGN8KBC3brEPG9/8R1OuGUSraHTVzPWP8e9IeVM
AOPRXvssYMpO2WA/1b9nS1E91zqdiXCsT4myRS57eVlY7sJ0OnP9AuOidQ+4dj/FEFY/YBLDC1Gj
2q0ylYh+L7PaPvoMXCLrPZZ7JUrDUSalx94iy/BQiqxbviUFEFWwr+VnJX8L462z50vMtKwlnTL/
5O9Kz9hTT4Bz4tCuB30g/+i8tWVQN6rUozWJYTGotqswP8P3qMha9q5u2MQkI8pjS0DscbeiG3iR
uEaJ3bLskqWXAebGzIIRFMWolkFQEOSpv3anZhWIwo0fGz4hiShk/EGrs+t5kzpy3KvZc51LthiL
yK6dHEo8sXoY6nGgk/Cf21igatqRjt3iAUk5dCDGamktHu9AOfw3K5eYuzAETDplqrJDvo6OFh3J
P2YrR+Yl4BvjKCp07zYcibxpFCzk9R31R06JObS4G2LFXIOMrzQE4k9iRw0Kl1J6GAMkKniQDIHY
L4Y1pz/KjAhSbQhtkTsWHkW009iwd9mM54rr7H6qtdGT2aQ5cPb5+O0qY+fPuD/rlJazRZH2eqbc
VVI7s/vFTBv8zTQigi97xJexe5Hf3rpgNSX2gZTRLqOLefDWMrYe6wMhvTKu2BYdQVvtpNNU0dAM
+yJsi65dik3Q9SkeNLA0NdEjSPDOT+mRKJeSLI95tvh+HH3S1dSoxxbluGTGCAtKedkbPDZtMGBp
ZLGJLcTVvFjtsm3Tk1EFsQVKUmnUaXa4KtzFO97a2m/k7BZ1FJgj1KRk2GGpkb+MdSnc0La3BUqb
XDL9/7NYiHLeTOrTm3Au2JvHSa3lAmTlYFG3vGfZr3L1sS/aQxpZoJyfbDubcrmg/tlcbShgJ5lu
aOAEZ83Sk4bjOpeLsexfJf81r96edjSMxWEzBOVrjdDAXOb+aDf85BICiNtQz0NJWK3yoAxcqnSP
YTN113v30fBIDl+yOeLZSJuEUwNFUJ165/mG6JwhZDyLvNow4bWZg4fWk6GZNSET1A42kh/B/v4H
OECQmfI/Gv9wEHJqLBryPKz2j9KAy9TZb8oHfgy6/NplnxKVlboI18gpcYupzlNGQ4eElcCc7wLO
64QjcsRvSx0noZnGQFWVN+c/gtmkm2S03/WSIA5bGKVXNsV5mpcwOY/rFf1jCE8SMvWpny/2BoDx
nZD+Xr+xEwEewO/Lr7zbr5mogOz1nmIPBgnpK1mMpfeKFReAPXUv9NXTO2a51Y/GVtyjjc4byJM0
vodgXPXN9cyzddRajs86ex3GxnqcYTlh7ajC6US1OyjCOGIkyNEZqQ7HU/rwhR7xRcKegQHcjhi/
e4OXWvm0BrvfF815DPCXUTdQg/2KyV3i2p6+elMYUPPeFY7d6MuRp8l0QXElpHV7LxaKbnVimRay
3R0gkRIlNpWNOO1ZKzI0BCRSnIiEh/AxKFsGLoWVg7lDxZYhzcssIk+HAgoQD1HFefqNwp+/I+Y8
f6OX5xl4hJeggFHLnQDyXZkGrPiZs5v5NuWXftZcgHfbkjWvUTis89sQh9v0XBihkmQ5eca/YlpN
syt+jcr+NbumGKAq45cc7FqUbWzK6S9aNfoUZQr1aAjK9xdG/QkDZJ6ZT59/93FYBKEWJfs3H0C8
0RJiaOmzi1h4ydWgzBu0ejYPm8phHE+q1Qw5jeSVDpWzF70VnU3C9soeatbERYs03pBMsPK0Q769
TkF0Xueaoo97W9gmkjfdRW5GdrdMzh2/REJpAZK+KmTKxBtywajba88d5VMhACQ91R6Llly3VPAE
aRvQxZ72W8n2eJfE3uGwFhUGmMaLXbuPVDGwuEJA+pAKNkhNTGbNt6GrD3kT2xVltafnek87w0fy
RpC7Bu3G44Ld0HmseUyZwSo8/76wp1XKbaK4wN/MCpiyTe74FhgQu1g0SUJX4H/8HWr9YHnePWuT
fM7ZyMBORjmI/6XGREoKU6IFKSICelkLSXjzRvjIhZBmj3ePci8NzyytsnZCLLVino2rivQKvL/i
3bKCzxFuYLuc6Q7hIr95S8Q9BwYqumf4cf4L36nbxWav4KyfVmZFmTtYKvxJNta2UsdG0GUtX9+R
hlf2GZBWxoU9uqzQjeR0TMwJq9KOX4xqV0z4Tiq4r/8CPILlIgKm9ldSqcLfaeaMaKmDxDwz+XVf
68Tm1ilbvnoKhyNdKb7uAOifwgYDzAs2dSCZf6nPu+a62pR2uf+EP6hFDv58iwhHgzZXe7rzF/X1
liugOSIbsoYDXLD9lZvUZxshkLkZzCE7DT5cC5r3wAd2ddkbmtvTCXfq87+W6kZZVUIJuQ5PNFpI
XPe6jP0hz8Kw3U7uWOP6H2O0rwnjkScX4uroXfTigFpzGNQgr/anZ7+TKUaLAo41xV+Yzkyqln49
Z5chO+sVwKMTbXkYmmjiA1laW6izHDuCCQYzn2A47ChySjfaB7GY4L+upT6EMDA6tfNqW+IRGGf6
B4Y3m5V3JmVjLUJVfgR6oiTqlidMySkwsu2BAMlyPMhzcxnBfrVS1zQm5n9kMsvuDPdDq0gU4Ys7
ZicNQ2JN+R75dd2+fMd2rAhvTFdAFDdl20gyS4Q8Ot9yPPjxvXFvAkQiHja+bc+p55OPmlZEiMxH
c3t1nEF813xfcuQQeR1BGdX49vUXWhC8qdHA21wb8D2dXsgxi60owFvaXjhcvMUf4V6cN/2P15TA
4LZccMXqMMaJruOjoG33GLKyjK6TPLetDymuPW16Gvgx50SArfWgmlYO9VVtoGU8kre4XI3vstxe
9vOXrPqD5MOnn2o+KoPN3Mqaq2rjKGbxNNQPQDddPsyzKnQ/dG63v/Z0yVOzL/qW/f0KpaCQiFjO
GBxTZJnaGF7VzYDKlOyS6QvYIXoZj3vKIQfYrLRwHFwjHQsd4gSFuauetVYpanpXL8F1p6z4QKAs
LzxpbAnJjyMssir709t09mpbyyQF24TJsdIVpiidfLLaHOmYSI1q18MAymllF/yi3hHL4cFbeDCp
f9qDQ8IUS3MU5PmcyK02Wqv1MEvte3eye573D1yKukx8yY/qtiU4qginG6ANifO0pbjSKTSpN6uG
amKr21kOPIJ8SI+vDxj/OFOmNtq23eKSUOy4h4jdERJiNgU3lP4HSvDFbxkF5JZ4W2qbc88ZR2ZV
Uj+LDzkab2X7V+pXcg6Ny8uTIZWzu/mUMOer27NRktnStwkIIB7XG1Qduv7UM9QV70Sld3+cJ9Pm
avHiNTvMZbg7/Q0fKKqPHhLgJA1iarnCjSTpLIyjnRGr7UgpFvu//q33cufF7GZITE4emUNXsMuJ
v57P2R1EKYHxCD+Y6XBfxR2o6fwZs8KTkDl5CRuEl+DZEXq2uLfhTFZd6hwGT3bbM9WMO8j9mx4H
9K57Atd/6kKRW2f2+DVp3nk0jwy3ejqRUOYChH+UcCl2bmTff+W4pVopVAVVhrS4YnKfi0QpNNjY
2J7o8YBX7oU/hwZbtw4jWEarLOGhFtE9U3QY+V8d0BiSq9TZ3cvhyv4fxSzCJcHAO+kM2uRXtwFA
4z5yrDSfkwCjO6QnAAqgb9GbEluEwuFfljr4xctJjHHwVIQ988L5epsA8SySQurC4Sd1ON2MQRiY
+F2XtBx5w42YTCVIvrTg6yZw8/bdy9WyRy2u1/jN7cqU+Qy2ueivXjKptkrxYiKLx26Pz/p/kLuZ
TdXjeNVljZYZcbL1kuNtuB7SEE6GOmUKZfoj5WB11c/uzAn7ZG4zVUoGpmkpPMl1xqUwe+U8KX0y
tKve5nzffk/Ylk3dUcyrql5A/44PCf2Cw5S5Dd0yzzpzgjtF6qjQtXR9hCpgoEkX0REmpQoVl416
3RMV2wQWoZl5mEm83eLG39Rz9hwqLx0WSicGpwFMrvsrRZB/Kb5Dnflc8Lw3MuYkA/oLFlEMPTP0
YzpxLRnMzXzZ+AsHDKuyADBY5nkqKkDwNjs3s2/ifGImCcn0RyRleA9Y1ghz7riMIGKxoMXKOZhQ
zATdLJRuySAup94llbxFIivlgueNAA18bJOmnzSUrMeIgn4jYFnYZwKGToxxfF/RP+Zl1KQazFUV
RSMclC69LQgbKKLqLWDRIcHLjVkDMxl3GzD6iBf2cmXn+DUmR30W+mnyjpgjPHTeYpHI6TRCjD1e
eP+H9ve+8QcHvCX08R9uj4lpz5eaOVaYj5agA92CB7SyxQmmJJ9LxBJOqyF/CWvNRwxR7lYzAXPs
kGnHnIxL1bHIuUICdHgN+W3NI/2hqTyTE8CQzRAsQgcLj/eJa/YFY427F0zy8ZJL2/9qu1gPwRQf
NcTdaYzUqBea+VamfsQL1Kve048EEPrSGvwWnyfZYfC/If6LIN1EkHLcqqMoJBo3jLCgkIdM5Qs6
kcLguIFp0hOSuZxOUPLSErV+LWweOFap2DlWKyj/o+d+QU8521dNBZQHz2RrYO8RYCzkQUPHximf
hI2twOh2y4zebRZu0LGPfJjM/SWRjJSS3On+YqlUxlw+898iZ91htRbQ+OMAT5xkh0dCw3IWpr3K
MU24eUmNFOv21Ow1fGKXEVGIBtAjH2hYB4J3JWEEH049VdJx9iOxkhiaOHx1EDQeksIiRgEDJpoN
TtgRMVMXU/6Iut8x2avPdjrybEQksN/PaIX4Ex9lxV1ZohulaHz0h0x40h3C5ux9bSuQ8seNBHko
obg8UThkm2O5uuz+oGP6+Pn85DE/tjwL/0GJAPPCRA8w3fhgol4Z7v8Rbr5+4WDS1qsfmw/kcwTG
SfitavsYbhIJ0xnyJ2tZzVTEL+q9MQDwT1afq/+ismA760vfFslcTdxGFvcXZp15/KEEXOigzZ+a
45w9iaoOrYnYxMEK0jhhnWcr0ieDWIGWZiSO+lleRxOAXOtvNijpeLvoSCeeSY/7OVsbt2zLXt4O
s7G7seLtR7QCgn0Xy3CaQRgPbc3XWKmH8eEGQHOt4AhxrXKOsK7myFdGgar1E0YB3CWpoSuiSheS
nhOndtCX+bVNkNbU+o+EVzgI0szuKLEGqklm7e4DzDWA96YrWLiZUBZvJ/KD6rscWVevjMxgeV/A
WrqN1gJgwUjzYxDcuBghfogBmvECWpcDmrIPAJTpAxpN797iI8ljQr3l/qSmaiOIDz/KItmN/k2t
H8u4bVWL87ujU6nYegDjVrbx5isMce3DVrcjrzGxZOUmU6K6/3Yh5nMNRmkPbM5XgbAzctC2gewU
mimH7NUltdCf3UMntbHgCA+06g55AMGZR0g325WosUMNG1lNfpzhPZufBiBCzN+qS0xopl9wJYQJ
4JxwV4knrSnY7CauXOr6ro+FSgR7m9+m4X1D/EBFCE+abJsxBCxCq+Ho1ZRcBe4CWdjgh4iRhmVK
PeqaVN5BBTfr1TezitEFmv/gZzor8T6Rm+ZZByZzamDjRlwXBZkRXKs3APR66kE/x1ChzdRO+i6O
WsOO5FcZlzNgqdXvHnS2ps5YLwTNDalHv2r0ac+DpjDE25ugpb2TWFk7a9cBsX5B8WAYTHOYS5Q2
5y/SM6coWOhGZ5s8WIth6xzekX936VstfT9mKQW+UTLyJ0nWBFQ2IySL1RLDeVrw6uGH6AbdibHD
poakMjwHxd8ZUVzpNcxlsFBEVrfo8umTTjo7NUPaRb2JxlIwRiEnzNRxcB8O5ldfjF7vBpk1aHNJ
BejzA9MN7axz53CO27cNIsNiWWHyvmGZ1SNz/RHFid2vH6Gha60itqqEjmgLf1XUbaxSmrsQlZNQ
oSPVhpv7U49oXUZeHsJOhlCNp1C6nm+B7wUSvSiRo/jh5ZQ9bOB4bfJResfe8eEptzlr++rpHY4/
RX7oMzF1+e7b943kZBwjGRqj+WdZKCU55aaRyAgcBQW074OvKlm0OsK+7NSAbcp0y4JbJ54MxOI/
GYhrBmKBlMo6yyz6am1uZmByUVB0nt1LdwI45Njds+sc03CtSrfxQrwQTJ60ah/MsZVEFfcc6xuo
SmNeC3j26RjAe58I+tB6jyW5tCCV0oTL8fR45TQGq6EGGGl0Dxn0W/Xcw5f+ncs/fn6VuLCTDXve
qbnXlI9f1tFFzppsLUhtOf16EhUQm0YTA5BVdVtnXFNPu07zEEF41oWIUPko9/V2xlmA7C9wBOAk
nsiYvOVWcpaml3kaBopr+seRLbJb7QCtmv7xvLrBc28Zok8VxSTnCp+2jEbXZRtVe3fssd1AVF37
bTJnZk1kUrOnW36hDBGyoU5mnBbCHy8ueJU3zoPruSd2fEvoXPrZW5RZqX157I3CQlojclmVOBG+
hsoexdFHYgFlut3KYjCyOiWlWpoRxXMYxAPVNP+AZlCEzfuDRBVq5E/YoraSxEfmGJFd+CtdsEpl
grf33v92xbsL/NXmOXYXtFKvJO7DRMR7SbF7Vc44M5OXQF1EikPW0tmL3Uq9bA+dRrYzu2h78/9D
rPyXidDLgzF6jxgttnE+WCkLQuv9n7aG3CZQ9M/4qGFgsyFr1/WVl/yPSglQKhpgJYTD7TVPnXnD
J0WZ6eqGMSlLuwySfLXMZ0RYpITjoSySPAdZLrM1KXv732z1dludFBIbUG60JYL+MWGmWeA2ihuZ
aCCjebcDMCrIxP833knsFms0Ze4RnAPgHMpkkaG5UXq6h1qJ+1Gq2NOotYOOyv1Kpvwv+HcQyF5g
iX+WD4J6SKnmtZe2U2OHzH6xGh6TmnM1Qig0+kxJGWqRewraxNPZgk554DFHDNMlu7fFuQwVyJk4
WYNWraq3vgVOyvd3NFp4FoWOjHe2dxt11vjG1JBQUFSsNqOJ14bFsZiknlNDCr+fXOHxNUf8VL3H
rh48yqBrLnrJxufqvkVQTqt4o9dFI20ZiW1HPOedLy0CQjLxe5rSBRSUu2OQKFRSFR4/O03i7zda
appa3KfwUt000zLXO4Us+U4g6H2KzRXHExc1ExZroDX8584N5R5U3O1gOjgO0sDbAx9lkGvzjuOD
AU7/CYmaqAEPdGf+i/es5ZnQQH1neDE574D63g0AktEW5i8YsbhHGBdAOI8K/dKpMcW1uNxLEbzT
veeFyrutibQmxleZ7UAZAc37AbJTMm8Pco94bBKnd8f5iaViMJ4HnGdLyp5PLAauRrPEiNw8UxIF
U5InJRT8e5xVEHS4rWwbElRgc1wDL6g3AqZA5/te3lUIjQ71QtmAJJL9yiY4j3h/kQLa5yHCPWwo
gcSuKP2NyUwfWbBrEBTLCHiJlM+TDhWEdtqVBKpUZtwJMbWRoLPeOTIDLNBCCl1V0eKb6vZZda91
zOaP6cCu1PdE019jcJHBjhtsN67PDuEoyKKWUNPaLRqx3p1oLQbDps5b66C4inu/f9dcJUNaoMqL
mR8iQ9tw+qK2sTzwzGMsuwn2N87voSw+i0vo9V0JIxcpXUyIQ4TyhyQOJdPe7RHOrCfrIaxExSKQ
rFrK5DCGXX6e/wohiYq0mU5edf3gu/J5F9+Gfc6TaMHT/sD4SZFtu+2ZQgwI8CF3E2756nR8klHG
HEiWffycqwHMJ/9jDp2uB245gJpNc9ymI0cIyakC6XI4FLlUMicBBem7ADovgJe5HDfiiEhWxScn
DC5yg5ALYvalkRtYWc6S5pvja0/omWdAkBZnIhw83RMaiYFtBTpLFCsOnpmtxiKSF1GgrOqdUjFG
Zf7eB+4ZPCPfWSAnRHD/lZL2A7rDhcbTjITEjOvF6F/2XFqINUBLEX7MGzToO/ODHlsQCftlXF43
IU3OooVd+Kkmx/FopwFyK4QVrr9C6DcuxMiwkeow5WYK/551bm1wsdf13qQqLvB8gvxDhe3vGh/Z
9jpAEIVGQwkafw2pKg5XyHxQomZzE4S3Y3q5prYUCWu+rMgMyAgvmhBglCipm1/GFmbE8YDtfd/+
s3bkDoOaLIQzfiypRW+FDvug5rdvs/S9xxMIrqjnJEIG/vnda6RJiFdh6OaLh5C19BrmNYKA4cMS
X1kNhd93AVxBifFFNwUPKeMLTLo1w931tYZFV8PnpGFyuofqlJ5vBDK4drtjHTdm/w/Z/nhbsuyS
l6OY3OX+j8LKDiU9gerZHSyFNbMKWTT3FQalFUkmyrwHoGPy3zj8+c2nlMgDhS6xa2ALg+/TwH7v
IASncoi6pY2oMbOmeR0+ZjezCEKj1IqgbBUhCuwHTaE8m6msUtiFzV+2vYCgylqUm64LC3HNiRbB
8pkTMG60vMd3DWQGGAYjHzu6te0V5fYdofTdrfJlJauITfFk2mfxtM7Zm45Unz3ONw7so9/bsJ9k
HCVP6pRyISCfAKZgbjNUeuppajTg5j93TUZlb0U5coYq2bx5gO3evDK8XbKJK7UZkhsDaFqn07Ug
1Ucuqhc6S+HJjRVhGWH+i7sWI998XdCrZ8fqekEhJL4iNDLE972RnXGvkJkwmIqoIV2lG8T/rKkb
kr8psBwXQhYbWpEoNGexRFqZ+7C2W8Z/wPIrGxKKGD0UjOFPF5LN4AXqcbEB+kKZORVo7OGuQ/+S
jWNFpWVGmqVc5+LTmF3ueBTM+kM+r4E2ibbFlw7PRGYT0NLpMxtLoQvhonMbUGA1t6TLqYRhNhVT
z4TEGtePOEpoCXHdZ3c7dFtP3qyTC/8p6LLpBlUQ6BNg2Y6HPl1polHrAA3rrGXbPUr9+avAO05p
RbuPXVcMPIFAwi0Z/JeKQpa4PKT/G1RdQYkbO0inPSiu2+7CjiJ+Y0bPzHUKQbj1zx7+y9F5MKmN
91zepvQr9QmLfdpdhvpNUl3vnVpq5pxeVt+CbzdThtnctuwBGBhNEmfRnyYZSrtrB0QTeXAaH9aY
OkHtZOoP+vdwm5T00JdfvJVjDQ516B4Jp8Ren+iKlZbmJ0J/EYlAb5FcrhMNGTtWU5FZZqeCJRtL
kUeqPx9uXIZPGwxP5VUgOZzJUlI9gP5x8O7l83FJ/iXaCkCGk+uoS6ScIzyoN7cyZr6530i7IA0v
ggNPz0rv9FTvhCnQWZttaW9psYjcE2N6j2rCHgVRkc/Mnx0p1NypX9njR2s1RdFgD2KWpn8BmJVP
WF0WkGVKxUWVjCGsEr7GKMqBeCTT8QjhTl5M+cxWO3V78TjoTCd/kZiH1S2qpnhbeOF7fTBsRfFC
ngdFYGUbctfrCSSXYCTWGvmqtmegcTaqljdAUF+ehrBUA2zaa8FzL/9zgS2FwXSkUuXLTyzOoUai
8887BPuq5aF0+n7iohW0+eDyBGPKxC3t6zz8MRl5DgIWfCF3GepXnozxgCeW5HCEic6ZgzVup+yf
crQ9E9hm5x1FJhZsQvAxkZA3e3XVlR07FX/2CPlqFAj0SK0xKAah7o1yMO+XaPiHKsxMpZh7LolA
Thqw9w7jtx2pY1kzHT0BjU2UpAI6tCOsdvYaIVczdwoo/MXoqLz91/9sr5+Wt2i0u5VsCWy2wuBC
84QwoSgVlu3/oJQY5UQJVLOuGrq9ATG4CA8I++yxcEb3KJ1AaKi5DCeRuYdrNUxzH/OeEapVdzDT
gdsdcAYUqhtLNVljfsTQmnpSon5R0BxlOYjB92fZcp3phMZQlJiFLk+9hG1D1pFrkBdIsyAlkg9j
jGmbVAwXfb97Xql6bt5YOM8aZxPDRDGj4hfEhj5dPvGV5YHh94+BxtfUjJt5uLBucpNoae86EyPl
343+ca9t+iVVgRkFYZbd2+4KCaT3vRj+qvX3Dki9ncfricvJafMGyM7eX/ONk7szo/5a59iCVh5x
IOn8MAqcnk/BVmmvS//RweT8bE1Ob6FnSDG0Hn+f77ZFM3a2GirdV6Ev6FN/etNLM3/4Ab+drKTZ
rDq3PhIrvHeRdtWbdBfEn4RoZCi/5GRJHZHueltiMaCkx4Y9nT3LcEpLmeNR7ep2IX/UAoDFaLn/
Exb5Y9Bstp75zT2FntbxBqTuPq25GBum8c2j63NAejE3H2x9k/KsuslCeylP7Y0wVERa1dO2z/sn
u5LFy7Wa5CLgWk8dlE+qgmgeu0SoT6APPpeYgr0ZFFLuvNuFFQJZqN8kBkRXUlqc+k91XOS06nq0
ay7G/P+T/S/UuiePb0chVp3eVLUppiUuPrYzup2BUVSS6KRvJaAIShmx0X2cXdw57B9UVpMlFUrW
5XB05RcEVohYAdskU7EN4SEiYHMqrr6juLFVDr7nfzN6ezxPV+siU3uv9MnXWIRWfGfNkmv0sNKF
+KQN0kW/iSFIcU9Bh7qiiD9Lp/1xHdcwCDcmCOVU6aR9IVKkudvCV7fymjBACtikFYsizU2Gm58d
Qnrjs3s2Cx8FSXkxud/O7S4lcy2CAaAjeqXpDH6iWq3nNXZYVtzq0Ny/ecK+R/olFo6R1aEYsQb5
txz6KNNZBlnYs0v6Syt80wloYJA6BCeFzsp8m6JMp4ba/zIAs+GopM6PFqRnHEyZPO7oFHYd/qFe
pfBbMBlh3jUE6WMeRfAa+Van2OPae4H+09oEJXr5jcFDEoasOQCa9+7rpKXfo4q3Pflo+i3ZCG+J
D5H60+HiyMsgrLWSrr7TP/L5dLOvFaz6jEGKmDHt6y7WJjDPnCvn2Zuky5Ybcdi+KUWfuSLjedeU
+sZ/U6/nVXHnqApn8c1pBf+5GSFevibXGVl6l5HqAGRjURXiyvoi6xN0JWMGadbQZ+QKci4o1XNa
/2JZxPYNIPDVLmxEX2z0NKHeaGAlC8GtyU5ifAbE52wHh4A9gLqX9jVUXHaBOtth92A1ZC1vjCC9
jQdOaj5oPVbOWPDW2lXiA+Y+s+3BNo4ZdSGvHXeIOHW4x2BLfamxp2hViESJ0sWIuCnTFdWPnEtG
6FxQCueFVJKmf+K3cZJQ3Abp4+IguFJ8k/A7DRnkTjdjfdv3AeLxmnZqDsGZqApR3cB5+YU7tYK/
B2iSSXC+bjY5Cshrt13BUrlJMHMn38szxDdtHA+Eorfo1hWiOsk/bAVGqg4/F2p7LFUwUY1UYgtg
UL0Uq2jVI2UrqaPR+ZJxUL5IKCA5eCiZ0xBuvWUG58vZLXVnj7de/th4VbWMt0I8zxV/y4mkovtz
Vzg6OtyireThp2OJB+uUN1B4CnEEUE4SGAk2I6v87bWdRVrbcW7C0axvxQIVunj2skA7wneMSOWu
TAgaPp9jmHiJLrM6T3nerx89v3+9OHc+1rz5HJlb+gE/r+S4vKOeP9VhJI+codpFXw7UdQAc62Sb
ojD2RxNnSq0wNnSDaLbLFoeF9pz4cVzuDvlEQumENP06l48MTouMgdHSPMiLJ+lJGa8zRQvrFdAQ
5+/dwAI2dCFJFXaMdoJQdgCLH1HLXPIqcuHdLr5+D4Z0vNcoNUELDYgW+XmTYgWOkLntd7o18FQJ
fXC3IADgrhvwJOGFqHG9v1dsUtpJPmn/JkQO0s4Qrdot6tsHAEx+wbfKw+rM70UD7FwDm3CYDw+Z
AOJkOKwSqvBSLs6o0U9zc2X8OTXqUbTBTvDWgClAoy0HNEHod2xqBW2prHLsqDstriwki3UGygWK
QH4E7bB/JpG+X9YwIe4KYv3kWLUzeGLgn15Rc34WuOzeyyDnZwwuJbuvBjNu8bl0Ye2B5c8Hmd3y
qTzY7TMXv3G/K+nrqEG7e9PzcrcmTPIZ95BpMB76ZW5M9ZLRk5PL9Q401qmoXwOPBomEEypRYepO
kZrtLqP5TCM0lGmHoUYieD4LpGe23b9Ek13CiW/zNQb+LD26ZVahnl5khkPEaZOApbxALS2/yVH+
avlKsTNQ5cg6y80BcL9+pyW3hSfmiRgd8DPx0XffM3iAHEAqi35QLupW8EnYeJppZB43t3ihqTWb
F9XZOTrJhtxKiFReGSp1pKdY4IYKsO0rVLrghaIRlc+ZUxLzjedXuBEp6CCTATfh3mEABE4APXj5
5YBlHUnFSE393y0pBqRoFzmSqB0KU4LGkgG359IfDXUKCdIitb+i5rdgvz5pGSyoKLmnoCDLgZjP
4qU1r5evOhF6ytM09pFwXTNLghZBcKwlAelu2dfhmDg4XfjkX/EdXQxUkib5IXEO3aaNcl+NNXsp
6nMkmZLusARdCSI1JDliYkgc6S+popHezK09EAZ8wAUKDwo7MR9iDZyMr6qj1c1qawmijwRFFvGl
QiTnHoahKwVJms3HWohTKOd+Q6MdqVU+cFM6wHG0fSt5520XIiJlHyZAAIHcbW9H3MtwwaCSvsPx
gGRo8kn4+lGMBETnEaFaWAfNMuwBTiMZvzpE2WNqM8sW5ypa6ffenSJ60bE87Euz8AnqafFRXAvZ
YbAaNSMkJwUoSUqryr+IMA8of1VhsoKEQJymFsStHoBO/iX4BcOum1NSNVpTu5pqivxakBsOqdot
xQx6BO6lk4J6EUyfhlMRF/q3jeT/AT7x8es5hswXP0z0hVAUuE5r453UnNOIjrm7MZW1tURJTPyD
G6wQd4jvQYlC8L4lMdS96y5Mls2bVzFdPhXfh595gQKwTLS/ZHr+m+urz1Buoxt7vbX5+zKNFdWp
pXg4OwH5e+9GCEBCsi5Beux8aW8N/m/APiTxtPij8bFiMJfRSoAh67LcNVhMs0PXM24mZl2hGyUz
FdpC864ka46VPftP35DMP2fDKYptweIG8b1LGsse/1mX/FESrJqor6D2UoBGjBZ0q/wS5ThYLCK0
Qw7NmCz7ob8AAihTM8LxEgZJwK7aaohehXnKE7wvWmOClWzUiUufYTUFEWq3RfeFESOocMRdd29A
o7N/hHjd4zCg9IDwnO43H+wf0A3SHA0fVkA9pTa71edG81wKSoxojsIZSFagvAyAgstzlM14+07B
YYzUDt9+btHURMhg94xP7GneYZlCVzaH2MQ1uYzmYZlwCWtH++YcXrT96bQfNZsQV+DEWejwDX9f
VW4E+Qz/uJR4AQWLaKnfbA52EWH1dZHZ8wChzpF4pmH2jfQxMUb3L6LIXPJBDeQIc9cvbYsRQVho
2//2IQ3V1IcWEB5QoPjkAcnvcwymtOuxR5R6M5MlN0xRKK4gK+c5N6pD0yG9upUyp7bPHknt9lBR
bmc3aLOVMCq3efvpTzBJAahnBhb+ySo/CtSaFFrQ3jARBvVMXxWiS3uKMIqtbGpBeNNblHwCY82d
z4ay6UlXhG3MVOU26IV0Stq2sluunKs3P8tnplqG+UZiGztM8Q4JusQiXSbzQk1Af1cov56QX76c
p1XQBL5B8UB7m0Rto6Y5shIDqD/oj3R2HyhWAxvY8ENzHOzLur12Vftee4Up1xV7GA5HFYpmDS2V
7YfybaHcP3U7QHFcF5QfIN6b9GfGAmNVxAzvgBpgA1AZ8IlTPeimLtJ1pCQJTVIZ5CHtE/M9JZyc
APnDTUB81Vm88Ry7ILHpFuyBqJnD3lpohGDaoKQIoh2hKlGZ7LbnZaf5Edhxbpzmis7y0AiEXtSU
//2ysQAg3W7Sr1Pz7EA4lcDjRw+Jmbk7XejqFZZyvq9XxNo+nhdJVyDdIq1C42XMzLb4Db7WthOd
3uy2jUfYSnaaZA+gv21ciIyEI1HO4X10qkrbKWa4btg5RBgaYqQZRxGCWKLY8JZZZr+dKFf8Ie6j
gvM6gNBtHrNnw7jLR/1MzeNQgilKNGikfbicWigzmp92y9Y+AGE1Tfl664jeq36cFu6fbu2Vn58e
PXjaQFMZ8X+FWS6gK92GdZild2Yf9HCwd5r35t74WTXmLe2Bl4fJrjdSD/6/3TqTZukbx5HWrJu7
fcmtodDoQ9TrpFKtfpdnH9WnJjnCh14JYFDSDKct/ya2ApK0GZ77UKmmkbHtDkx/fQnWeAZ/ezsW
gyX+xOgUeIE6DDJ26Spb2DschbIu+cdqsH2NbuY0CWesbCKqYsdtu6/cAbkhNvkAxHLfPmGgwd+i
UFnf9EeU469cqSEr0lxf2mxRJ2VEvPKnIwma+9TtpTL1PnkMfBoDi/HFSC4hkMWuYWhSMtKElHUZ
U+KyRPhV3gj8Z9IQmC3h+XsityKuTfhZ5CijQNAZozr3qTcUNsaI97x7L6FsEmwUy5oFYBir8g6l
Qcq7S77dLc+z1FWz/M1hZyeWXHuV9AZMoHzGSa291LeOjZI8OjXyeRlGNX325TriPdANBQQ7EAmp
/jOMKUcECpxAI34C5tcj3Ke9HqQf2X0Ba5Yn7wSolF0L4zJBWoI/CHAtq8Iznaan+WTdJq9fKLDh
/fqJPwIOZpCUsS3Lp64zfAlia82V1x+NsqJEhFAR/wE9nrxto4ZCXYcoCpoUv/E073Yrwr48GCJY
eGBKy14e8osmXb4egYKt8n1SztaMdzHJ9bQfWWiY8MBXXeGZmOV07+pOblGqCo7IB3beiAdibN2c
/YrghjISKgNB0DizWgudyJFQRMNk4lXO/rNbDvA6VzZMx354gcHHa2EI6/Hf5Me5qJSGiG2JFUCI
DkfMAsroqlkeF82T16DaDeiuSmX/Ha2SEE97joOm6maJkcaxLf1dbeWRtekavPhkDqJXnETztkIh
oNe8AV9B+lqBPaZYAcXlpQkHFMRoTnW7EL7r8tT4L8uj0AZJ+lQEdrXvqYwpJI14cBUHDBC+kVFD
3aIJAGfqXJIikrFyJ4VFndlcbKOsO+NXEKKL9iTrTOxMSC+WOu/sxYtWmUTjyvFRuxUhgtq/WfzX
r55zgoA7WsY9r/jODqJ3ghK2ZuCm26Sz1d9AISCKH2Y8YQgCh61L6i6wJTyep8TP0cERn7KmyIm3
8HXz+dsRfssTaVTyvGeLi0hBbEGdIWIsh2VM23WgXLH8+CBXuozZPdUW42AQulRri/vOHNi++NXZ
WQOFK+uaZ1wRSf0DKma9/aSm+2R1dmuyvN7x8sUbx8P9m4mrnfdE6cg+1f3XOxliaSs7i5ObmWRt
jmW8AEzQZrjvIN3mgyK7KP1mE/OmNXr6oX0Z+sIhoRL78GIbPVRz/3KzKqqcOmNJEJsm8q1TLL7h
vOrs2Ud4cx/e4ipRtagjCZtkYW40Z9smddj7NFIrqgaAtPhuafn72XKzK31w4SYt/vm4fFQM31dP
a63KHhsK6OQTplawtzcnWGs30VYpnBJBoey53FKz64O2HIn81+Udkv2TK5ZO0QSmvBOA4cqA45gj
y2Q+VutMebQG4QtcW0ktk+sOd9gtu3n9vOgdHJwLTWWxVhBh2KIhmhUQgEhOKJzML8kUbR5crpc6
FMgW3fyDI284iSTfktBwwaGUCA63n1ZCOxnNsx3TlPwBWUP1/SI/sIyKHKHWDcejWjvMUmBWxpWK
6CGb6mb5loSfBHSyBzwAqz1rZ86LyPQXvTeaqdZjqgyCGWYanZzFfNzk0dbRp89okbsQ7QlIwCpq
inmxIVCHphjIAHP8I08l80fj4Nd8M/wZ+qlO8Ine4sW3eQr3YV1gy27vun/sAh706OoH9gGiqNUg
XXAJS9n2pOn+t+ueQ3xPqLwmChikABSqrx1C66V268beL7ZmGMVaSz1I8zpbC2n/d1IhIRjxOZiS
itctQPWyk7GRn24+D9faaLR3vL5UokLVlOcWQ6ANsWNm+NLcnIPqGMaayv0YlaWmHdNxnznI0CZg
6apAAedaK9x84fyl3pfFtqsm2BwyRqBnkDiI4J+B9LHRd5MH54ftT4C8W88aVZ54GA3UACxV0pWg
hYNW4dSqXyl8JIlqRUNzBnDu3kz4r35+F61JENXdxbsnN012IVGRIqlvGAD32DR15qSzXAYzMwXq
u+vO+IQN4plU3Mw9d1RYu/l7ScIO1e27mn4vuzkr8Cdp32/bBx9Smykqu0c0+PxE5RoNUkSnyqQ/
Cwbq2RHKfJfjzYYNTXTxStiJ1ZA9E2QAv4dPw+17hV3KE8rDr+dnlpFio7rG59ANilDAPg6FHrSb
VRyYYhVDP/2d6Qm52ggVta4WThCsltDRPkVnEM0r9wyJXexvRrydFBT5Kyl14r/oeYv47BSXxj1Q
Z9QitGe5/Xecs+/GpJFIkHrSpLG0R7Xbrw9QGtXyO8ZxgFaOXxVrP9XjNjqvNZ4TKqyVQbr8XPCI
9n+eU3f/1o9coibMK7XjDRXpoFjABZwHqDLScdg9EG1q8SZA77pDFjDuGXcAkFGJFeBhpQclt5O8
b9L4sYKcZMxpPNn6cU4kI3Ujl+QVy6HOaYat3voxzVeEw4POGayUiLDzmGfYCLZBRWy9fIkEL8e8
QraA7OjlWYksInZdFQF45pgVJZ7RwODDaIVzR3FhmLr3jKRaNN9vrqdFulDyTi5UWomrl4fZh3LG
yVtRLAEnLDevg6Ie+vB2z8RyutikNq7tMaIaKnVanngVapVnjE3RiE2jAf/LG6cJadYGvvwKI+Lr
rqsbBC56s9kj281hLayI+utWpk99zDX2eMehvLP53IVv82JxmJ0VNYD1Q2lBtn3Qf+NnjFyYRUWl
WPJ0p3/4o9YPSXtfNv43UZnjM8tmVBReqa4ORqCGVIVfRd4Rdm2zS0PUb5idM2tqZMCnF+aOxR7G
pkMn9bu1JYxoKlpRaBoOW/O8Pwhwv0hkorNX6fS5g2p2tuuFGJiP8SS32AipPftYO/Fwyzk3rGGS
jOFdOEO6wUK6AcgKNZ1D3ERKn19uUYCQmomLRw1c8Wt+0YV3OeaW6XQ7yKT0hWa7b7HMM3nqb/mw
jOPYlW7btj27F5dJOKmwaeG+x5vC5wACyuWf0nmYPrCKF3MnoBAojpguOQf992LwQX4rDl9vtmws
hZgXmPetA5rxdUrSbUnkb3FtibXUrDnB4eqGccs9qGNDaasnl/pcpUdBKrfWw2mogq6LF+wnoVGH
uWGyYcYh+PnvsyW3JLAkA34XjbH15LYnw+gPoYBJ2Zdl3etsnpIrSFNvjUaSQFFwt4rD7c7fAHLp
w0wCNJjrtuenENiphxjFx4oHSU0/TarM7a9AAxoMeued4bevCtl9Ss/+epZpoS85YnqRNHAYYMpm
GkDNu0J3CmGb5BaF2JPqlvipCoXYPHAfjy6sVki5a7miipRPpjEIfs2B0GLzCWi9DWoZ9xgGkLkC
64MJwrFRXMO5kQO/oxdSX6sxlH7VTR7JtB2Rqr8ZZsSfQfisomErlAfW5ViRSeqd9msPn6Dcgp0m
pC35tnIjylr1CpfZ9+dfPJPFMD2zUPQRiG+fvpV7ZMGf6zmYe/m9iDm3WpucRJIL1BogPAnfqd/3
GVDIiqbnN5FO/MXO+zNE+Jrxo/rW6YTH9cNwlkTQWbFbQYIneVb3Xx0pDLGkMKlkTgTH73g9k5gU
gkOtb6Bq6EkUpaWBLyXYQcwQJ6m49s9FuMRkdFRXaZSCuh8y7fejjCYG2CrTLJu7+clb7yvhNc1Z
OEyucVQ0Yjss1m4Wx0o84o0hdJs4OoSflhjao4CI6wvBV6bOerSt+mb3NCq66OKUspZ49ac3Ha9t
bC3qWcjjOgFXz9evU3ENiAxIrOSJBSqyxUGN2H0cnoQ/8Ys1405TlfOcz7Eiu+P3zYIwnal0k5Pe
JsYrIq5xCVI2NKsAI1TTVz40QtcECi4h8vMv4o9ERH2mwCqDGuu7rLbGPv4mgy15geor0ndYeKUG
Nw0xQdSveVWPCrHXvPbgP+23NE4j14RLXfw6CC0GXSpv+TMfW6AZ0kTNpebKEQNbDUMXVHi7Fp5+
1RiFehys2EWL/Xmt+TWMvxG0vokK/LeWhuWUOus0A6jKm/pdqwwsP5dv7A9QZ4DK9eWGlJOz1LeC
sDlkiAItFfzJH1/MvsFpeJJpWjUtJxNykcJ8AM2kpfbMEBf3V7A7zYzLhEw3xpTP1Qe8O7ZXhs29
Ud2283FAfnWBFd6tqNMoYXq5OrAZW+r2jUpdmyoBsbElbIjflKT1ZYtYauomvX9YM6jvR+H5kL7L
jNN2aOXAde7y2h1nN0U+snNBmmKM3BZMpu+CP91nqVBAEoauS5koHtl3j93J1YJ0iKJuHUD+ht+y
czL0D5nq1YFszaTe5hZESQk7EWc4UulziWzq5VHT0xStZEaRkTuS1gTVUMLEJTUeZql65u6o8Usi
dns0vzXeGeXEyU3+f8+ler62Dg85n7nvXutA1k9NC/Fiz8zF4UJzlr9/B5WiAs/wMyLa5MSFjA9F
Piivztm1dM9f83jeaLKIbLNo5Xxofw2LO2LmX/Kyw5zK8nWkq9HrJWYT8UCdHab+za8n/inSa88B
k4cqq8pB+5nPrT4J2TTHQU0X92eaBXaBriNSMpG1bLKFpGFqNIx0iHiZUwAKg+srbQqFrsV6GAMJ
QK7YEzbMZkP5ED/RpmaArdYFcRdB+cR0ohT8f3yM5gaI9vnwpb5Pgjk0mI5PxNwlECH94aypT8zY
OprBVuTAS+9uFqufBVb8N3/Bz0p9sGQrBeiwn0y5zPVz8sinAJjGNgqHiiSOMIXS1y81A+OLA7Uo
xdVXyEhePqQmontrZhZ2/fZ/lG4a4twIffNw1Lh6mXOHHNN6WAuo6Uj8U8s7yarA2jOqOutBojUq
4C5qkmQEv69B4z+XeIaJkbUZBCeRXgfkY9nN/uYSkrZNCLgfKG53A+N0MnPwCU40FWTAQ0heE7Lj
tr9i5vRqGZDPmLyQwsYJEv+HpnTKrMG/2TkkN84/YGZFmtLbtj8x9idxFNIDWDFd6WpgYyKRC5QW
0sTKEEeFJ33F5xMfUR5EAM4sCNwcsS0btj1n+3e45v7RQXfo5T1SPjoQQ4D2J2HTAkg2wYmqU2G1
tzVrxY4zRLPc9kJK9q45cR2Lmiy1B7vIu1nBSAFO9AmiKIhXv9YrBd+U/IdXIZXrDFqz5rpD2chn
LEJVRtKE1gJ6Mb1ctR2Qpb3WOwHEaz/kcKdR0cWX/zFuPIdiEx6/Cg3GB2BdkU4vau0cNzTDA8S/
RCwOTgQUVmO8DLS4Cw3lveG6VRVGCpmKE6tRed7PCcU/kdN1nwJCVAJKavJRWx60MJo3c5a+tmzm
QFjQCoac+r8u1xWo9xAPZ8PszG8nUQimkMG924qchWglfhBNY9hm3YYvcuImmXeoxkDjqHYBDNpp
rzQYB8ErDTrcRK57QDAXdApUazqVF0WZFKOrCW/FzoiQi2ntl/Ht6beWvwhcA/U7l47qy0w2QTrq
LdrsmVXlcCwhW1mRqzfgfsmh+9DQ59bDyuvhYhKQWh8kL2F0l1AWhVbnQgJBBLU4pFJz3VUJm0G7
SV4jUVeV6AJTazWKnOqVdT8TfDyZFEi7hOVxLxopfh3WSAM4l9NYhGZ6KoEXEcRr0AKwS1GU66Dq
IW38Spxz75n+PmN0k4KtobuH1SCanxtZC/Ra1AmtEerYVMz4BuwB6mkRxTk1tjx63a2YMvn0rP6l
nhTmAXLre+6as84kZ7PovMUxr/yJMJdP+g9aUuCt9lCpOIl3ax/+kthZPSqyBoSES74Kl0HfKEwK
ISQ4bKhnBqfurEON8kdvJjmb8riy8dtqBQgw7jfVCZzZUCT/Bbh3YbnOKmtTIta6bZ23Fgzfw3I1
NU7dF6rxcAkUZ3X4KWo/7zAB1iTThHHDC/hiPQ/3GaZcraFBMVkWiWcghNQ8bagLNaWmXQ3ejtYE
D10iubPXZtCMks7GL3+s1KxvIe+Jmv2+ZTgaexqIaROvEfau7cPWgFJJNiiZMRJbsNyMyR/JXT9s
rDLFjCCsm4bsN7Jr8/085DazMQ+yy5iSWM2tK72KXJc6gx4j6mg+QoTB7Ir7ZI3BIe44qP+npp1r
qBrFdM5HMQ52+2UzGNbDVAjK6EJ+uRJW4POyivSZzUeQq3iNlkJc51aEvzg/yBc/ozc9WQNvWtCv
6PpqEX/VTX91yAB2uYmXAXOWBLzydR7Ni74n7fbg03EZNAkPXSfL1ZIs8R8HhteRdjpek9WuLNhN
8hnJr+n7ItM+absbWEkKx01e3xU0CG+Jlt2sY+kaPxmE1mfDilUVqHIGxdwcGi6rj9e9cTcWSyj8
A9PzIOm8JavqusH2TrceTUw2z5qgk39nzFIbXCY5ueKav2xG74E17zzApUvXmdqtmB/awvvJ0Mzn
6dGF2LxN8UoAKsPPFwUrO9293wmeauxfriRpjEcbHxVjJWRf3WoHVUwJT9DUMRbI3ZnSSlAKqpcH
pnMgHs8r7lZl2CwqPyvNz2wYtWTD9tCc14noyRay74CppVzVTrPB1syiF7h95CTDFl+ZJWrJ6PDA
D4opBn2qpSdKzyZygRbpeoJluA4wimeoQLlWKwb+oXCkwWtDMvKi/eMK7Yn6nc+8fE7F0ZSmKQmA
5vUA/fbh8+ztMkxib1u53qV7jySCOtcQJq76X9+eD4/rF42fEYXCmsnn8U9HtESBOCofpn79ZakR
q210Oj8pNAcxZs/DrVxpczO2y7oHQ1Rf5AulSrIWMmW5nVMfnL/8WhPDDMO7IcPfoe4Fv37dEBU4
DhvInDn1rlb7V6fmuRPItgnXsch8YB/x0ZyBzXm9ra2XwbgNb9zFQNf0sxDauoTZ2czseu78ZmLc
WEOFeK/9hDOebkiu8h89f++GjVpjO+1T5edkIz3YDRqvcX76MMVtNO7M4svyF39QbMMCdIevaEcI
VasQzcKqkT7x5BV2JPBL96HeAJMFKWBrLZc89uxmxdlQwLMBC7qApy0m6hW2L8Hk0/xGCMAVlctb
6Dq6wGO6XN5Cp/AEH6nQACJRs3ww8U4I+rffS4h6cYFRW+UKQ0RaUNCz34q5+PoUT4g2Q3ohLPHU
AUqrh8Ntm8/tLM2LmryPIj8ijjFjPAwrRhYezrKSW5qA1i5CjaIzLu0Bxv3ordtJVUO+1H8PMQRw
2IYmwmDDLQYU5Wxg/w8WhH9EtwL800UlmsS7IW9yGuIwaSB7ztGPJ5AL7lrPtJmwRKxo481Dak9/
y+3V273rMpYCNWeCYIHuPYziHdBXHTzs36nbA/oQjlwogn/0rXIZ1CzAdgjIahfYGK4IfrfgeR06
GYGIuY+kQXsYkFsgirZklIFhfyA9cpu4vCNT1lqG8ypy96WYBxXrux6+kI6atKOlyVqs9kslQTgY
qkptauh8j5pe2C2/VSw7eAGydNeb7sfzpQG+u9bmMWUOH/D5mu8DbrE3T4ppK3Jy7dDM1kp6RjTc
ydUN5UyTPfPoYOQ0vtjySKWxhj5+9tMjbNAq9q3C/+E4+KFUn1MBWP9DdZaIbAHwW30TNO6Z5AOn
JSTJ5STbjK8ZSVCLmoMbGbqJ3JjkBfUbYodSdyWafyoH9GijiiskyK081e7FYbj1wExwC+B4PAKP
rhTjvQFmgSbjvv5+NpR2p8eXdakjMyzZ+vFBvfFGhxj/R+RVhxtKOJJKUqkaqWQ4JOnN6U9RUq17
wZYzJtPoQhP48xYSArFq4AaplyFvONPh1DhtwFIWr8xfDlNLwSikd82Iy4YRzou+QA1pn+nGCypy
IlgqWB7AGlxVUCP9q1lLbTX+I2io1xrufBekkQJlqpaRR2dZPnolqkUX+s7qT1x5W2dZCCtlUMVw
peaHGXBadcYhjs95PZ3cjFlcE89mudJeQ41oAFwcvNct3MjKjSHd6FW3LWp2/J+EKDtzGvpEoTto
7SouK52vhS4LVDNGZBq8/o3Q1ssf2YQMn9GYgBOVQZxEPkEdkTJYdcEjIPS45Z5DHBpGh9dYfPUM
9YzpFDO74UKLAcYZOmRjImWGksADx6o/vLyoq0IKNIZHpzerTXQFxhjpmYyLF7gRZHJ0qp3ZoYPf
xa9CNnPf7ol7X+opa27przWkzK5ETEnxqvSTqGxkn78hKorZTyg896p5uN16Tz3BGnH63zc40Vtj
yDEXE1UTOpfV41c5aLOGYRfSycguoVOUTquGQuaT0sRDdexDl0Gl131Poy900i40hdEMD4ES5Q/t
lL+2vlubdFSvINk9H4pbQl0msOp0dVj2co4rXtPX/2s696yDBbC95tibDeEgT0w6GvqZknXaArXo
yXnnYc3ikSeTq9NMdWPlXS0sAZ2ejkGxUFXWQGPK8bFujdrN1ZsYL4OAsSNFqZdkwZexFfxSxoL8
o9QFN71ZhKaEqdElnMQX+mZG/zkBSNs7gdRs7qNjgEJXY2sNUNQolfYA6zBOXzlQJzrS14QKWDoU
4vvQ9XM0HplT3/UH5+xXULtvHL4F85qrw6Ez42zUpf/bipCkhjzYjtgcmgXDwU+fZC16nfAsiJj9
hUyC9yXfB32P0ATSt9qA6KHiSNZn3aJPfAjfFBXZDyy4JPmysxnCgJMjTts0Nqswg6ye9oPXBqF/
AapLaMiuV1pWzK93RgjaccrCXuSEqLmJL6n8hBYtBn14IzAxcQVszV5q2ctlICwTOTKVIv1fhv3V
2+ivjGB+AzOri1Gb2GQU4sdnsPFyp5HhRaXmAZ4oyKhrZKH/KohTxxMl+cnWv1iKN97w+AJpPtwi
PAyWUHU9Laq9HtkNRnRJ6155nb1kpIegE2tp8tqZSvziyxDW/CPj9ZxbQUtQZEXZ6z1wNxP50ode
L+vB4GJZ0t/HrDzJ0fN+6usqGCkjAXZ/IEHQDQTR6nW4XgfIlVcio5BLOe/uQxDuCdxcNrH4Jypk
fIhSeGKK30FS/XsgINnpnxBO53Mp5ZW+vZqWgjWL/QkcI3d6Br5bqW05V4XCtWXdG72+neIpY1d7
Ujl7hVWYwVqfD5hDVwggaJWBiq1qxZVzS2dthT3cbJ7oSbYK9jUMb4H5F96WD/gR2VqaAJSqJLNR
B+pOXRqHYOPwiAFj66OcDqPGOlRct78FEeTukQm38aquqpwaYAAhkVSWlCbpeTHK5vDA61XkwPLH
AOEDEp3LBZhpZRnwa9M5jg62GhjQkev04HFrEQphlgCmmiuP1a4sRbGMxi4XaQQiAsLmDfcfHL7B
hclcW86P/a1GIiG7Pm8f+1fa04I7XK6DxhQ9/FijJGxD2a5fWNH7uqFlGXvXxTOvUd8PSTqrVj5M
J5Tj65yjowBRHANC0pAy1ItAqi9pbY7NZrJLIm+0Prqb6/Rx3B7U76BM7XcQXyM6ajolotkGWXut
jEWIVPnHxaat1MLuV4pmGjO5d5kQDld5Z6vfJG22h4oLctiORvCQtoU0ELH4v+MJOOpVVWw5bo3J
/zEprYbGpEt437CpIwWoW1C+3Sc/OH7f3PTW2DjSqEWyldosUPPuhAz98v2Hn7d1//LAGdSmySVt
1X71BTbM7hMaZd/Aa78YbOVQHJ25o7w33wrMKCvaw+hqb5qtFrJNRUfLyVAtUmenohIXJQUjaDfp
Pc6a+BlPzs7r7ihXoKmFmk6LW4QtpQ0LNq+rEPyfUhuJiVEp9BtiYiPC3S/2itDOL0bOEDbCqMgE
uD1hZv5n/UXFlwOLi0fUbP+xhEG9IcWySp3IIwLLCnQBr6VjjeoZ3BRUsKJT3NhTtj4bzgMniETA
Lu9EfJZ7IBu90YRAPUHwD9ysQsnSxQLu9Tts2CvaLb1WkmCn0hFga5Xrh2+pGHKj7DhUND+21k5h
+KTkBgyqljHs/RlYANsMCioEPGdaWNKJ2Q+Q7+NJLlMXnwlVvwtD2OknQ9grMhhK0WoAtzV4o/34
p6jZjf0U1cCQ2ehBNGIsrXY3E0/SH0FVkU732HEavNRud7XIZnixd6WCbBaSOCx8T18f2d0yl2N1
s/TL1pjZzqjfmHIhJhT9a52D4yT+PYKzVz79Yq3TDkISJtOaqU89sQD360HW6j4jQLQgaB09fE44
Bx4SObdtR06k9SQDD9JKrOnDJiA/pWdFHggchpq6Ze1TTbRKbA3OrHL+fAxvEc8wcmqbLNfLZjcm
0ZbDCq8Y/Ph7/b13XQVAfVECzF3X2nApzBBzS/y+5pngJ8yrrsbUEMU9jqeAkidv2qqt9hH2FxuE
Or87tIsPNtWKFZ1YHmfhAiBRf8qS7098C4jJtK+/YN4fzgKu+IkfsQXA3vK/JtlAdXFnhgsyP7DA
eQz3oCM4F8eu0YTbOWwzH1S51vqkR1jD9HcrxBhEnTQBddEAen+TLdnnzVgW12AObk36FzEuncL8
O4VBEF+7ejNoOq2qM0/myxdURaNuxfHKEz5HHJcdpXmiU6FajkRLh20ghq+Pf+d0cRPXDL0A98J9
JTaXp0v/yvuAiURnRmGv0CxMANNS//CDNvYDgmT79NqnvIDKYQHqPTrwBOcX0AHyFVTWli271IBK
S+D9JGC4sGtilnlIkvUHIDhvCx4R4ACMc1TcnDuhx8uEL+noMB0Vqd/LDRipPSkCZxmjN+UBCbBq
c7fIZLVCwrEcRmR5SoGtPFEr1dUP8X+9IHX8E+3r2JItMpraZ1EjFWXsGgTvGyUYad70T4L84ui6
rvIPtGVoQxxq7cwvRzio0129Pg49O2aLQTPrjGyMmC9XFqbxIlmETGpjl94N2naRl7fPzNahajXd
A0JvMPhtZMyeqOwi9ntslx7PMFvNkZTepC9BYNBTEOmh4h+oqLVcNXnrQuVlIPrJfpc1gHYWu95+
nFQaJPpZJIUbtJBFlQ9/wawxtGcOf4EVEbIGgk9Do6K8JnK7nMgRox4MRZ47FhDo4s5eadqwt8b9
8TVKwzTUQBLcSUllk6xGFvm9bmV49/xqQ+E25eg4F4rCOyh7s+IVMbqe8fiVG8doPi1H1hW1Taf/
mZgX8ap/w7MtvIVmpVlvIKyi3YxNclqRCztUusY3bMQesZ0NvfOuWhvhyiGSOIqQ/lSjEPN3RXJH
bgV40XZjVBsV1v22v1AW1370HL8Ej16odc/8hTvPtkSy7eeBTJ8gEPrHcnnyOXGncxGlD3CKf+Fu
96hGFP6++FUbas9PqOLzxE4u9rKHg9TuW9j1BbpzEH5rnRfyXwkWJXZnFdi0PNo7dKMuo5QfWtST
hoIi1tG3YMqQ0PIHLnVn8/h4KIROBZi6t+6PNB1LTdmCAJioth2SBOQAok310pcN5DIRwc0PKuzC
imsAGcFTPbukJ/bDbc/cRAIL3ED+UoKIYe8IpcCSDYcJLosinaAQVsP1RNRgzh8uXbC/l4BXvdTY
PodDsHfqL7d/2iGKbb5hHW0zzchhRV7uYADE+0/bp+iqHmAnXLYAUI7tH7G2tQ6Wi4USDqjqoqV6
enVTruWjca3j35KssIsvLt0MiWC4uujTVVHeENR3DqWdD6dlUNol7630KhDchqJUAFENd5b/hyfY
J0njErtBCTR8CSMSL/0IEknNQwGOZDtptFYkP8w2Wwtum9buKOIxvDs4qlOCZV77YL2Bn+ACxHTc
OQFyAfVy7LHnzaFV+aE92whOOIlz8AAfe7uAkyjfL3pHhr30VZHxYztbk8RsZAithxjBDEGMY8Ma
kmNVM+xi63S7GRtDaRK8b2ivwLtN1PG2MrmUKExhNDCP//RZQtPxTrTm22e3A7J5jJT93otk/upR
jd3R/TJ4gtIgIAgImWe+OrkObND2G6VJKVq9T2e1LPAW/xzvEPXsXNGba+7+VCqVyDCCxNOs+3uq
DdQAv/IZ/2Dcuo0ePcl0rngCKKb4xIA2rjKYOsHCBiKfuu1SPcwXHvw1QyREff6+aokzte0IcC2X
0UWWJVpdXOwWtQ+MW0WWaNqzrbOwqZRQcI+6xJkDLgbRH2h7Fslb9j7F5nk+5pspEnLXPmPw0CjN
qRtNaamwainK6R9LEqCqyKtXJVTlD2+cu8OqD2HPBJbS2nhvo61H4bug9btSFw1nQGoCcsPeEK36
3eXzzPuw/x0FT+2c/OACs9Z9XG8tCS6v4joM+/WbgJnrtUhoshTO6HZMAiGI85SrOi785dR5m34t
3Q2M45LlTJ/1huhFXfcLGXZ4v26G/4HEaV+zzUoDsNp37OONUZkvGPHc3IJAHn+andECUZWRLszo
hNaeSBs/LWUxZWa/x9QOZZSiIp/yEP7LBBLxUM+1V9BVeNduCPr+j5jb/EmA3FHOss0Qsckv22ey
ab0Q75EXoXCwQnMlXpsWfAbE04+Kq95hFsJGeLGwJ7qX3uxpI9l0ert4HXuOwSn8spuoBtbdQy+S
eXp6vbxH3U4B4370jqTlebUbruOzyNhwq3z5YJsVMT39pUhda9Eha2NEXnQLCT0wsdesqrYFlwS4
0M8UW9suQ6LG+tqsa6RvzwdTbXpHiemhvw3VCjQTg8dj09iI2Qi7js1RdYqLz5bOfGIRdi49ZZd9
agd7fO1Rv3MBvw2exNQTjJASEeQP2CQJpXd3kCJdHOM3XDi3acO2deQW4AkieEoto83fYYey6YNL
ePSQyfVQUamlhla/JbWXc2oW7xgEG1Ey4L4jky9EaQ6bH4nsYfbXFGKeM1xIMKyJLtkYit6cZAuw
jWEG0Ku7uVV3XGpQTCFTHBLlMy9RxqqUm3Pev6AsWEALKP38OsD5lsiR2IR6PXJ7OeAXoG4ecYlf
YjJb6WUJHrPCSWeY3sQrUq1aB5+tRW83vo0+wdilA5veqPP97j436sJ7vXFL6XPNxNG0jhdDz6W5
t9msoKQM0ZSct++/IJcaOQURDN7aDFtp7B+jryulMPO3x6KL055YNDfXnsogsjy6gzVspsj5qxi5
pHGsaEPT0bSxyRLV+sjAvs/47AvwBtwrJYFCS/M36TzUg5zAAeMr0eErw8Upb3/fNoY3JZFgpG9e
8/CvEaerinL2ADzrkFX+IUSHVHuSltOe7Y/QtmpwWk7xtwmVN5xkr6BY7U51uCpKZVXCgZbkWaTz
qllZ2Jj1RgINTopevNXoninzvKUPcNFlJc2zpJBrS2cbTj1KnZgpb5D3blyksbGrpoq0AwhrLyse
8ZYv2v3tSrbbmgiCUHvXSV7ECTlXZLiQG1TbN02xfdodVZdv4e3QeZ7UyGvnr4yHBYGYEqHWx8N5
SFcaeYl4M/TBtMWAVU+5Q4iXA5JrROaWOvrDTunhHubZ502XWPly9iQ3iiRFa61RGoy1y/jqvfV8
RJQF455QcQDAxqAGRuliK96B0OmzkZSKZRZJBQ8ZMXwmV8suRo9gpG1Te1rygjg5Fg5+jgd4wTXf
P7zIU+N6H3ZDfWYBIUyDnRIyxETr2w+uUSdMfIs8HwF1sx1Hbm8YiwnxL/sFlXzv1I6+XFqPM3jf
/MOL3HuAmU4le+xQDAag88d6md4DHkY7bcsWaXMBYcSb/AabWPSsflPVPxzYpshyPVzls9aMqnqR
6uIOJarDaKVIHfKMZQDmfY3U8mMq9NP8f+1QTIuIq0RKFmThBS3PNn7DgCbkIbQJamFQ+ptq4YVW
opf9TovaNrONPnseNKRYhsNafEKOVoNyVoAk9T1iW3curlEDUxMvyuo8jSwon/BWgkawilcai4JR
Uoz3/PNcyRJz/02GTAp2pk81DPQ7khzOPNp1+4tc+pHcjlI5DhbGYw3kuYswyQTiqTKT2hQMABro
oTWoQaEod+HtGO8EF7+4S58QhDk4Owyab8RsigPxPZMpXUstyaKGaancio7cIJ8u1yEwv9z3tms+
hSumlE////HfujBrmEydawuJmn9NDqKW20mQZKC6m76Y3EihXZ57RFmeggZZdp96kFlvq9nXRR/K
sJ6zA10cmQ2VMz156ul1wojNXxmQzGdh1JsoNEzekmKmtL07oocY+R/wbmIPXOVplmiHYyCD8n/+
GOJpS3SUy0+iVO2jOxDkOCI0kmcVh7IfRPlzHAGLerRBrVj+36VoNxSw8U7yRqL3zaEzaELMsW3s
q5YJWe34PcQ7NYFjY4CujZAQ+jwYA+rl7GaU84YC8ZE71tDbYg/cTqVOME2LPudJQUJa80553KCo
997gKdgPDhE0aRgayqSh+y4EUf2ukJzOku5MMVpSMTUiOn4EwWLG92j6vKMhtCG4pCHuSPwDtFDn
1OXspSpMoh4+b8kKVzqRrw1cigODb7ThRsoT5XLLcZPNFO1obwSiMI3ivnN2qyXiaWDI6XRxzK4U
pINZEfo8SG8rr/EJDWy5phptbizNYOysDV6+4iQr+7QVH473ocQafIEUOmvTYoR8WbEE7clKdnTj
VUvGsfOAP03T9rV+AWX41BWW0geOnC/eSBZRPSuE/I7KpkIlrRvBCTaojQpQVf1qYp6ctG/q/lDO
EoelaTRTvS3Tgs38/UYy2jVpXZekpU5jtsUajPQb974s9eBR0GjzMYJk1etR1DMBMWxNT5dBReij
NTbxoQpaM73RmwPVYCVUMuv46WWX/Qy3dnzASOSYIpvDra8tMYoDk2D0kRRsB64gIHQ9AnY+xGGU
ByTL3WDztP9QvAu2uPqfnK+3Zm/Qd3XOA3Vi22DOKRY6LzsF1ieXAh+VrArQTVwqwnCItbeNOF1K
7Huruv2yWyUaLtfEZZkVhJ5JwONJFC/FddmCy5Nkp7Lb/38LO6tQ/9T7rAFF27Aj/qLfrJpu69BH
FOjyami7DZidMZLO+yZKeZrbWEQfuUTYvagz7IiGtknD64qR5cJAm5tWGP/31UFJUuJn8e7LMoxM
IiBRzFrgU9hXwLwUqZNpAJWktwvWf9OdPfAvlSanJ4WSaH4Jd935nFSDeTWJVzEGUHiBHu2rL95g
/XoF0f2LYCm4mw1nQ9tvzyMFmF/bFC6h0w/0qkJniqXSe88PNuWmTVJkRJVztx4H4Jy2RpOwSsuY
EUnDQFCje7tMddMLvW/rDqpOONx0Stia9HMBwLJqqOqKdtFIhYXjnRb4+Wzo2OgCExQ8Nqj70DEB
EcSOki61ID7j+RF4c5ZbExgKQVMccyqaD4EwD8UNXc7ysjAZVNyZ5xWMiy/F4a9hZ04UVAsN9k1/
C1QuNr7h547Elez3uYVPKUG4reEQed1lGO9HLleAICwfDYc+C+sz1OAcJJ6jgXgjE7i24LMK0+qx
NEc4vURSAcLRX2Wht50CbOo357Kbt5tWvLhjkTa+L66BZ1JmAuO7sIQyliQaJ9kSBu5EfWAX1tTX
IJoWsPs6rbMZC60T0+c/L1GsioyI7Y90YzrcyYiIqidq2QpebDMfSxz12HmAsF0vErNfGXonmy5D
mYMONDmDAtLtcowGRSW+LmLBcDfm7zrP4jZuzStyZInd3Dkp1uX9/z0rWWE/BXLtGo4mI+3/iwq/
xsQPvf2ZAVfy68w7hCg0Rka379tQebxlrIvL2HK2xaVf8nV7S4BmCsLPcLukWfPZv3wL9pvTw1ME
gfwhln8ehf14L0qDJ2UphKPka8JDtVTzt5UveS7Y7L1vzMBS2nPAfuPBDwMhYLA9/ngnEGlpPO7+
7I94RmKEIZkNVQAM2Mx4egmTMclfZFuyoHalhi/tHSh5+MHT2fceb7i9TzzJNC23ajGCXcX3rgzx
2kCa9eK51jOjYfQtz9oQ7vk+w2o9/HSjTTJVBeGEI/Nbw1nU72ctWb7HkvshleztkoDe4lFUrcXV
E0+ddxw0me+1NxUyIfxfzV/7WQO9gEEHvoN4zViWHKtnhzRBcFT5RZ+a2XkrKjFs26MDPV8tm5pW
BDxLHBr+ZTsme32GIznCYl+zxAkPN+GQK/dVlKUdrCVnJN/2Yk6wYRAWs6r03auMINsKLxawPpin
sxoW/gyi+6YYA4PtReZNf8zSnxxVNQZRGaekhX8YINgIRyvef7ORYWJy3ZvfBVKUmbrhpIfk/ABV
7rTGd2O6F7xUeR0SYXKFQcW4CO3E7Rj8wdot4h28ZbH0hnAuUOM6K/0+URbsegzseWDL7KSeQhaj
aScz553RqAzmnczZQ27/ivWEgs+SOGs14tKycUNMGIOMTFXRQx0J9DW/JuLAs/lcp1l5+e/m5zVD
V5U0h512HREiVP39Kc+ZY0ZH0dXl2CBaxIUsmH3t2BXmYB9cDgwpXUGv2OmmTa35iScLOdHy2X7D
t/qdR6f4dK+2tJUPk6pq09ASJVUUl3BsgPiDia08EuLJX6xK4XG8PmrKhtlVRHeGLZycsHCM0EeP
pWszV7GHsFTFLPjOnRbZhN9y3dYXDlPYT68Zdm8O2eVPggVxFY7Q6HbS/w6MVifU0gNNIulzmdeP
nPU4aZGdgssX/dlLY7HM7B0tZ4dOx2Md4ZZw/K+rGQceNRPjsms6cdcWTE1PMCKcm3+6fUHMWnMx
Ppfmv0r11JvDscK0H0dExyJILGgPY4ctTAVTJIHjwnM5uqSiJ/gyd8jgzd60COpeaq5nmvNz0u6U
t1bC2/Bhu3iIjfSZc8CJzuVIvT8MwHpQMOvKn38cC4G1MhsklyPAM3ADXO7+jnBKcaomISA5Y7Z7
doYW0/MbEW+TsdTJSrb30wQrwzBuu4LRs8M/Jj5GbWPIcEOb/rQfyEHWZLro26LQbWGvI91YCkmA
ciK1ehFcIpcFYI4hdd4Pbb+S3yAEN3LzVEIiFXb5GAZQ5dGP3siRDPoceJZkqBmNwOQnsPJQOPQb
I18lliyAI62BDROex8rRf1/uoue2VMptB/0rPR6ywnSN7Y2Khrs+HpRVhg1CztULSD/XjufV3eIe
TnXc/rMevNREgttwcppAjFEPW86RoIT9gPS1tQvJ9tCGfHhvJkWxYFY4YhXUa7f/31LcmVxIJBs9
V+KFHbpCCEjlPGy/mNa7W8HYfKEWDRIRv0nTVISXOEBhwIDAmE1Xf0N7PuKRPS0vPrJBsRWRFYBr
s/fhZXkgtb9XKJYqPys4G5VovTx/kKfr06K0xizQc7x7qxRY60mqMAnK8R9mO0BvVQ+hh3PPxsoU
dXXz6OdriOchR6Wb6XGM3h8N+C30I//yUV/XXkrUSsmjTKUcaFjVRMlB0E6YTu7tyrTuOCND6Qsj
DP6TfBnK5KsF/9t0C6BhawweVk4foGqlMyktiL7BVCr1RbSLD98mf5Vgsskp3Dk8ozxUAuROZ27Y
rCcUjj/U1AhVkY/zneoctl3Jyd09Qf6angJVGcLIEw1Dnkf2AUQEDs+aTHQsoEqGzsZvZJO15fB/
rHKXqfRAAS2Wxe0U0A8DoDxB674z5SVq7ag8d94YBY7Ci3kkeadIRJ+tajM3inuqtOaGeYky4gXx
01J/JTfLCwE5KeGb2tO+1aw7NC3EvmuM8qcEhvhYadLmsx6l+EP1J4Yl5uNEdFQiK8d9sQvsXwI6
fdaZG3x/gt6eoVoLhOiIU/rAUwVyfrWw7oWty2zwajVHWMByVFNZK4/UPkDxhbfIihjgsV8Mnk/6
tsDoP64zpcnz2P2p7mZoAHqq52rtXrPF2LToODHnJp09wV2f/HOzJ2AezbXNKdpXsXPvu43h+0xk
7/JVS0aZUoHASIJuQ+72umyFFjyxXBqFuNfFJLmAQ5SXXfvyANR7JPbqtevm8Gj8IWX8FWl/RqWJ
YjHBpAouoZp01yDUrZHTHW2asJGch0P4PQ+aCeYMv0w1291MHXi3GbhpdRTf0W5UAr/MhxE8ZR9W
8L7bBPkBftmWW6M31fiiKMQ3QPWWLjgyMW4E0LOsBJmbBul/DXKJctPALxhdld0cUozqFL1FBXJn
BSnCnDbnF05S/9YNXlnGIUqBEVr/AtZPdk+g2bMx/vG0E/fxhOsI+HcZKCfM6lddHUpcHHMJfdU4
STYt6swRokrb4C3GOMUfpeBZNCGzqaJGbXjzCMR4d15UhkAn4juI5zWLow1lvEyeqGtTfLpZZm3l
LnQFIM2r5wbJY5szT7jqZcUBC0qeBBPETsR6KvpVWbacyKn0OjKRgw/ePozI7ygFJ939KZ8hmXaN
lT3ZLGbM0cKpt4zUNznfi+DebEQen7JzWBmwe/Z8nFXomUCWGbcBCdEBYCW32ZCqbNmNgCgsjcoQ
Ls2NPRyKR28K9ny0XSB8Wuov+IXymapAFq5SjWbMiwimKa/VDPq9FSbnGfZDC+ST0SCFXYu0hbAn
dTAP7D6ATSQcH8TNy1+Js8qaiX2WAQcjMpk1D0HvTzoStn7Rpd0+MMitfAvuLzbgqg6UMlNoXqZ9
5CIe93WdIakbDuR3AAvBYO3bo2h/yVfS+pWUatVCHZdhUBLB2JHZyqRUBFaYILQoW2/QGQusWfED
GBRcA2Y9vS9uJqGNwulF9gEADi5eh1G30Hz8dLGOPrs7HIFzaKUnMM430mTYSxVczoos/jrvBm58
yEpLwDchadRIRfFXbTPzTX2eB4nbeptYYntvLILiSZMMM4EtyQMRTMufTp0pw5jao2A9iPa9u84p
VuSnIwYaasMf95pc6Ub7hwso9eA4/S18VFy1yEkgjDPhY/Ju2GHLPL+SLuYlOJ0E9zxNwMXaB87p
j+2CzUlFdAvOwH6GMMzO5anTE2vd+Xgg2DNBou6qvhY+ia9HNFk9nYqsV/hCdLMmjcTqoMvo7mxc
yileU0qdSRNgDyzlv7b3WebRgHtBY+4AgN8zFX5GUWNemca1sZTuLUZ/Pu84r2X80x19LPGIuaI2
kBWE6Pv1VbkWLSnMhJ5nlXCaH+hNyQly0/cVpR6cF09BiAEI7mw689T6Tp+kAKQXsg0m1vvO2wfZ
M0GQSgy9aiOUQWRndqSle5iRM+xShOQhqlbQ726BhpOu//j+PrRnWTHRtnLsfaBQb69dCTd98eEP
c62l37HdYWc3NDJYgx28da5eW2O2I2in6n1KUa+edmfM+MDboHbKple4BvzX8mn12gO1l1B+/kKX
PQFidFpjnRdI0qLfLxhNMZE/Wvstr4kl/WMeF1cRTQxJQTbh8sGj71WeoyaOiiOjKUEJvouzd4tv
0gqIuOEyjNm2d9O+N30Df6pnlqC2xWloBU0qBh+C/tnQfSCCE8vkPLEWpey03viGLZZCW8EUBMJX
Vgpkq7eDgxAm4xZ3UR8j/P/MpZs6jksv4uJ8IKlrc6g4CvKPqRF9r+n/7PTlvfzZ6WoxkmpqDm4A
M4y1zDcygNhhW3JL95QzypviV/vXdgon/IIwhcDLNzailL//Ve+hJQGOk2OKRmd88IYf2Wefv6bt
Q3tJ0tKrnoLIH4QewmHDPRaKsCRssltOr8RkboEjZLgu+qDYuKJuiEtsaUCrOcvd86KUlFpS0i2B
WpEP7gJF9MslrdOtaZqfDgNze2pK8t1fxYBqhTxb3YX9dUF5aslVqeSRZiMH+eZPWr1L9yS/fUWa
ZKM2Gsp/5YGRhXWSnk9RKN49wDnCWM3bHOHnKUNesU4LL9upffsf9lk/9miDmvkgz6nmX96z6hA2
euQltGaB6G5F28AR4JsK3ECo5tS43/d1QIs0Rf3ec/om7+Gz7fp5pB9oPPWfd1Ke4F0lv89M6j+U
no3Rt8CrQpGMNDUQUVTefUq3pZg44hCHXR/+jLLh/RK3GI+U5UuLc/vRFDGuS0V2UWFQOLvnMuVp
5yQzB4RLAzZyh8EBbyMIfEQew4YUzDvx7J1RZY8gQeeJwXPOqbPojnpcRV0WoBzii2ioDPWke0ti
VkXISPx+hE4hhPZFznrFI+jwvwRm9Fl9R1rl8YoZ3I1I6FOZGsTKh2GiT27yPre2/dlx3jDxXxtj
vdMaM3dhBgHIOvPf8yF/JwoVx3fRMOplAKouLa9it0SUk4X2YWmZsGVNJG/499T78+CnohtTNs7G
N2Hhxp70n7RNECBKSFl5j+9rLbmkjB0SgEQqnODSxwauWiu/LckqB89nD95uSAbPuBBbqrcWnIol
foUqbS8yNPgkfJzVkdfqpLrSB8JAmwbbgbaqFk1E+EJRwApagsBA4fnK0qsm2GnY34xzzEwSySKz
RLfvR6c27GSeIc5a+FsJxqPf58lh8c1P8EgLFHzOvHkS+i+4WveRANOtT4+rZP3brxDJ5NRRKJ8P
dYuOY5XNBqVq54E6VY83D8acs7ZAIjO+1yQvCbVp5Gp+kXgERubaYXQjN0aRnK+KqWueysXLDF7v
molucKTGkoFoYa67vNCcFhzDy3o1Z4XfsYvcxTBYvqnKG59imzL7kBl2sxIKJeDmVN+WiryvGqvV
Kp7myHDzojzKidVSnxVO0xckAz1OERlsolIzQNDSiM31g7xbVC+D7ncS0nhY4w2QfIK45McyFBvU
YC0J2tY2mkiklYnEBFiUqgNjLbwXdyxgridoQVeWxgt14PGeRE5hbz3RcMEQqQP9n8AJRLO9oJ89
AyUle27NDcrJ8gb94IGnxz7rOeiw4jtIYoj7yyv1/0OQTTBrFdjkeZzqvfECK+uqnI/YRB8P6cpk
f9rylGMwlGPOS4TIOwj2frC6SAvJL79NzgRUSzgYNmHmuNGI39atHOqmtPLsDGE0x+t0+RfO1p+O
GB8YPW/hdtHtcRr1U4RSctASigqLlbDsBH/U4r9nSACg5xMoX7pkKXUX0/1UqnxUMfWDASis9YPc
dK4CBbZlVbUKlBlJharNJ1K44HHbVaWRWKyCWPJxxaqgA4YjR56b88ua47uPWJEQQekqArciw7dx
BhiA2UM4ZV5OHRjnuPjXlsXBBr+E4+cPLToBRpFpld0Wk5gQYge6xs3+O65C+VVsVdSLy3WlfLTt
P7CorS5gCYEckctzPeQcrF0GW4JIX9LnWSwxxKbWQ0HMKwK2vRSd+tbgtiLiyOrUNHwOF+Y4jr1F
LmAm7OnuaIn8ILBmcsPFTdGlzpwvvHwrQ2De81amwnaF/YOasOmdASAPwjTa6/KNp3rXZCGCCIio
fJmr/3Lf94Lu9zl0wxBQ6qjgj791ygLU2vG1tf+HOFlGPRtbUTitHRiAKZLrdIznt6k28MupTtt/
/5Nt0/tQ2VG3B2DWI7lStiCe7mML4rMILTRdkh2GtuCrz1TulKeHPUAfkkpDfl2wz2Vs5M51G87e
EpQNhdPqyLjm4TOHTsq9aA0YcTIuniXEtD0quRVJ1hMNT4dk/lPbrxUyGSxJaOVpu90Hqk5zPMFg
odvcZPfTXpgdY35pNmsmx3LIQoQ25rcIRk3VSEFUICI6ubukCQyAGhamdsjdauufNFM7wXNYFc08
8wO0fn4rchY66iVAfZuGEiEzDAarj55lKMnodRhz0OUEWfJshkyXEZEmSOLFaqkTWG/+Fd80tcf1
9WOCiTuWLTzTkxA+q//TsPn+Sm3nuDHod9rauFgPOlvU66+hgE3X5O0/To96c/GjnvHok5asGaCx
YGaMMusHdkgRWgDxWe67sk7FOKmHN71ArhomupcrLPeQaE3rnMXYrnAIIN+2MP/uNvhW+BBJ39Z2
uGviqnVnw4xtcNtJAQH/nLamvP8g+/07tpuBeTgnmpjxqwZGZFvV3s2q+3JeKrsrLCzMtt2SXCKt
YLf/K/7nXuOq6MJPkq4s2/U81aDUfUdpkoOrW/i2jzlDD9ip8Du6bTadsdp6LjVoeZjaQdFuZJQh
qkGAfxtI5lobpn3uaNmEb3DjKXfMVY4NOhUwLyvISR06R2Yg7Bzhr19pK8pKvN4BghJrIxIftaVY
yxBU1250gmgzwJadmFnuB+U8/1rAZLACaK+aaHK/aU1WhuIfmT+N1bW49DG5enOEw1ll9kpRvObB
9+8ZmPhaqGICezLpQzjSE3DwMwIrs1MtgLn1e6QyrnjgzZ8nRMdDDynbuNu2RK+B3Lkq6Eif43Co
1hZjXgsVYfVEY9q1IUNKeIUKwQYbk3TBt8hYoNkQyXFzj5TrKIPU1brJuK3zOot2YsyLn6UcdlgB
xZ0JUEyOTbtS4yzXmx3aw+IrHADi2wSo2btguuRv9vogeCE5LCsESuCBciSUDLKQMq59KUTQA029
lDPnoZF3KBQtfSAFvYn/baQJ2Vyu2rC8Rlaa65/tr5EqVu/Kz8md7e6T/4Hep1KAMrQ4fWRZAIb+
PtNsn20/WqouQ/HaIJv7luv/F6oU98I8ShYvmHFc8djP08zcH9LGfkUEYQ1R9cwIe0drH/JFhhqy
Bb6ldIhyZ9Os0pEBS4VDLMe86DdOBeNiyY/ZCPvqPZk/uMkuCJ07AD9b5n+pAr/mcaAkbMKJqR69
N6VjEaB/vOtuQP3Gmd3WMOYaZ7yGU0t8mZgCuFtAyzILDEUodv2IRibt9RNeKR7bw9WAULEqIi3C
+92R8fuA/DVYIl+s/ykvpg5CEev00WRCSH5Ul9OygEO8lnGzopwmuwHdug/aWZ/xQvMU2WTWiQiD
29XbaTe6gPXELy4Uc6rbKsEQXuA3WN2mWzKuI9jJhIlxsMOa9Oh9kllIIQYqWzAvTjzeBy9+BIn2
XBQ58YZL/1YaugadYqC3PSCLPe2OSdBlq48VihDptzcZ3pKHpxuzgOJyppbLZN+RJnKyUI9H+FRh
K2j/8z13/wBUCDGWU/lPNxQwWbZLmjre6G7YvvNxNg4KSG0hyUgTds5ScHWzBsEup2ECjdRq+1Ua
bHAEsH4npSiorPFAucx0f6oTa1sqnsgEirq4LEV5z8tnsFUQJcKjz6PSRe40EBU2d/b/TmguWV/F
tggj4NqGjhgwGkrWTqGI0o9O89AABtsuN+P01o+6Xfo98o6BRYQmGD9Mo6K6NpANesc2Mc1oyhlB
GLP0AiL2M3iOHE+TODalHcIXqbwFE6M1cvRX0pPD3KMxWgWevoeu/zX5FiDnK9zP+FraRnjXNIyq
FR3WZHb2xQb6w6qq8GtPg7up0CjL7e0+xIh7zsAk455oVPFWCPbAgkX0Iy2EzQ+U5mFJ02uBewNa
zgKgR2PZmXcttq/rX6kwtaXcOg/s6wY/pQJbfPGCN8UFCJHZ6i6jNOkIZzzfBVqvrdyga9TnmO0s
qMhtWUxPY7njFGdAX/LZA/XE4BK5HFnNUUkiLeuWT+DGX8p5n5vt90b3v19lXxyHYRs1QMN/kHXB
x8rtpbmA15R5RShYxzySCtlYAWEgAhMpjZAfr9Yc3q+b4Ce28J2JCMezfV2UVN08azQj3WzHsvBe
psQeRCyb3Tv8aFSfRt9mKER/JXA5F4qSJ4Y2WYnHF7+oj6xBV2MkwTJJgOlo3UsUY9XOeECwzKtN
ItTeoLnNwVFOqqtVRaXL6GdNc3NtAsgTUrEJrDZD40y9IyRjKC6DJz0mJcV/z//DqMGce5XuDaN/
hU2cDMIj0fNenA8c4JuVBt35PwGfPphM3j98PZP7ldi1WTVKGscwGkFpOk6cUz6lxkm69Z8AkxRI
vefPjzitkXLsJqbOsabIqqFUUNyS55WhX090qPK9cPh+rpF/8a6E652dRjAETNGKy8jSfOsLjTVE
mxq/Qfxq1VxnwylWwwzs5Jf63GpfSCAyYmpJ/PYrliKUrgKY5kRpSeZ62xYbKycbG12h9GCnzOXz
3sGsIBKKn+S2+WcZzs1K+jhDDWQcArZeN4FifHbMn5Mqlk1az8QQgtUa0AxQj8a3fn9PTFWA9LA6
Rmnpx5jMKikS4z4Jt4gbww+DvzF92ovI7yzhFXu6G+lJHxbBCOCb6OoedgL6JcY0kaFut9C4vwtt
XHcVx//Bq3Ps6WHWsalYcGojXCPiDCvSHjrIAev+uAqdrUMAAS8xlS74PK7uHW7fqFbK/eVT3j/9
xh/78zD7XIk0Ki9p2nzckPbFafFmye0f0g20HrnOSzhVdzZuUBfzrZ6J8RwXWnvfI7iJ2GDprIuo
+ynxuJl5+eJ/FK3qmwjwEfNJHDWUluyXKDu8hZhnDPMwUceXfI0TO2UlkiNrOUAJtnZ7FV/33nuC
FJy74gzM1sMjaPEhFxNt09qeBxz3WndrmCWXAGGJerAY7tc9pjaC+9zkAZgF5KlDGVbzaOjG4fPn
lpGxENRP5vnmBhn8YpVsGIN0qMjZgJqS2xLk1GxSSuvJsOsDOMdrra4xX8KrT9tw8c53LHH3bgKQ
xTqA6pRewY0ANevtzMMyrdx/l2imrKz8ccys/t/s8G5m3kUwqLFWSjHJ3PPy2e//eJRLIeSycVe+
zvEK2PnkRCSrNBEN6Rogq5tiZV4YsEzB7VBVpaKQrQJva9Nnxa6M4EV+pua3RFGxB2L1dYzqQ12i
Lp4ATRCBmdK8gA3yFuDdc3NcjKYTmZiv45Go/BHd8peoq5GyesnrlHbOBTJ2FXjiDHtIPqabnG0v
DpD/UNMlhUn7hTey/lPf5HeXz2IUaRIyvGV8VMWpS8BhApC2vLHSrQaDsXSfrRASwDBVbgfidd6a
BaMNxaNMR6oNqKwYtl/YLSupNH+Em/NSpPOeRuTL09E6Zhk6mHwkunGySnic225gyyfH9uvmH9/D
GPu6U3VUp2DG+M5LEX1SdAKLGpVkC5YOXhzNIf3Xy7fN/9ui9XJqxyB73yssAmHHgTUBOJKRvfel
+oMhpcVVLm6IxEU4DKXib+QmXuNJmAv8HwNX9R7GmWYtQH5CuqAP22f6kq7lIVd/cu2f8Bg6TqPu
Z+HDE8U7cXXW64ge8tCsA6gjc67Bi3x7eUj5V+bog9VDro0nxazPeEy6u9QsQLywd7Lk/h0QDHM/
bWwYzOCR3kRu2kJnuvRLgyQn3blaLNXRQlmRLm/jxsih/5q+N1lgCmIXBiylGt3KCjguuYCeGfdo
NSuTRjhAJykCZWQjykpaHgxQPj9VuG7mE9hHk79wcshoOoH0B/cOAsdvFCFWty45KPrz9mhrENX+
8odRE2m3iIHOKJqt1DsKCeGkQiyvpnqF/6uosHVkGoc6/BfkOqgnLZ3atTA3br5zYkqHnI4pdrjd
VsjmN+zt88ObqdgLT/J48tJBKiM0+cBZyCdneyYuvFhZL/DqdXAMOrUKK9QQ0mhwwuu5dgk+vYKK
NWjbzMvS9xvqkvJnWno9B/iDPc/nnkI0Oqwxmc4zXHKBreLgBYMtMi6sZAraBsS8y4IccPAiU1Db
9bCnNI/2+sIGejhhyZuHeXPOzWawm8HJpXb/mcHpFQrRwruhlfd4qn5ncME3PAP/4wyXYzsyCmRE
NjD0y0wHx7kRAi1o9Cgi/QM2imR+MIpEq1faybfiX5fNIAy/TaHtBuHAzPieRhhhrmeRiin+OWFS
Ub3UCKYcrUz0ySgsOCrV4Lrf+S5umUPF3VYq3S4pEL+UId8vsmKTH/SZvrxGySPxC5GNGBGCDyOt
YH8f2ytZtW2xGZYoRGL3L3yhoGMoNHWHl9oR35GFgbI+5QA+Rt63Lm6Eujb5slFzmEPs7wh1DvLP
xzWtuq0iBOOJu9KJGJ2kfaEpwBrgVWQzdtgw7BQK9I/ZOChmwTrbnDL+r1KkNo3aXeUXa2AFDtI8
5DEaAbwLS75fdS1HzsdYyZ3qvDgQqLJPvmWf0VL4CPfdaCVX/p1AWpqPLfKuuG6tdwsWczvDLYIc
vupJiqaelWWk3rMqaZhhqjS+uUzfMRfUt3QOvLojGelPZanzDYbwanyjKzo+jfrrUbgV5lfJJbVf
5FgyGst4f6JN96W5ZR6e5/CX77/W6kMLlZ+mTcpjR6VNWR8ZkjxjaX4NEOYQt53xQytp1J1qrym3
r/n4SHBSLRwjj4eAFkSCOYOEsLZXa/+EnRU/TrI56CX0EaHwTndulZWKFx0ynnIo9uVdpvNljL1v
9uBSSpqYRs70vkQfOvx6TsGB4QSwbQbr8mewyS40hymbPWWpIIcfgMCvRp7S4AE/4C4CYuz7+ehr
ZvcbLJLtQSBtj1eAfp0rS55AmfToZpszqd9yXAtE1rzyl1vmltqarWvSfRp8aUJbwnZ2H60NH3UG
TRdXJQaJufC1H71ym8UaCYOpnooQVUSSELkSQeIDIN8Tr2GNNRU6jVY+xiuf0T6PnmYU1K6/L9en
wdviKBCHzGhJ70FTzNK7NVua6ouuSj0xK+rLYTzpMl35RmevkKcYj/QEIkcSCfTL1ngqqhewUXBy
A3N+RSNYGmTbnasolaYC9PKcuNdTPN7cFxyZHznnfZwlcgCjgMirUFb01qw9VDoDlRMy1ITv+3ir
Zg4+e6DKGXUhrW1O8+pztGoRkPTB14xcXyIULBtKGeBJIH0YvyTqAO/OchJREv6AH4hyR7HJalzB
4bnWZW+APr0sivxzNb5eaerLsumceCZVkaMchDf72Z8CwukzHfIM1gB2Q2dlA13VYFTAz5+6MCid
OLC42ZJnUSCZ6gmiC9O1vahXIe6w7lYAP+C5tUBqzWJJhk1ppSKbt2qMcUgeRSUhHWftzzqrNyfy
D3PUveQHwWwCUK1Sls2BD7CLLCe04JRs6eWCPU4tgcRBxDfXT+W/rkcwUJEWcLoNNCCgxOJ6Zy3v
pfP9hapMyT5jIQjlXYy7EWVQoQqyyvxrnZwT0b4ZYRBltqSpn61zM4JrdBCtpF806c3BOsSn1Jpe
X3/8sJBr7YlSTFf00cG/pN80jydFJEdgOXcqWfEMe2Hhb+vWBtmqLOKL/F3CspF3jr5FpEay+yKc
rX4UKpB/SlbkpWQrVfr2ljeVLnm8er2A31QbmrlhyQxB7CWlwG0ntB1E4oL8Jz+oTtBpkg4cnIYL
rAFZO0TQ4aGNEG4zzExxt/UVcCsooUz8/gqmvkJQK1veKBGk0zSDpYEo0/vPCQfhcWafdSofMG7x
Q54LUgV5Qzoj6rmsf1YrYSk/qO/wnvlKW2s7YNbIMobD3o5D2lFlsU3lWeIhGCqIzh7gJN46viAy
WsF+1JSQMnzCcyg3iqDx7qEF3/YXQUnz/uaN85L3sG1haravtBt2xJJeJdhLLpPxq3aJN05CeG7w
4G1Jl2C2WP8KzZhpB23pf7PDUm8hwwuCG5r0Vg4uG2vYhaL0p2fSqgsUvaK7kmjNB4/0F4uzjsi9
G+jpiSUpaIAFAcMw9ugUJgYX+hb3ZZHfx/spjYSbFRw/SK63dw/a7Z/pq2Uyfk8IMtLQD+ssU4iN
lfhRisQPIv9yJUt1ojN4mfTnvlp5tkBY4bNr7FseGnqtf1LMpoIEcclxCBSCI7/hDvVgd9cnmmaS
pO/yCcKRNKCYZ8w97G9IL8FlfvWP209rrGx3PRpEEhy1WdJ8chW+sYx8Otbcro9fI9Q5IgIboF4x
5XuEiVGQCn9AZ5zALAShDCrRSxlItfmzVCZHO/KcvWFzPZc0IPTO+4z7y/gWIzqXfgDDpY/I65s8
dyzEAeFk3sLADZfxy93NC/nq+HOtqep3kAkS+duEXFemI0ihhiKBftyva1DvqszG03VsfYGCL4BF
UkT6Cw5S6HH2/8O7+uwQNVa+ibVablb72jsJaEbNKcdgvMr+HsVVscWTP3axL3eAbJrbj2zTrn7s
sP2xiyvpjpagLYhioye7wUtaQRbIh2T1xxydENh8I7sxNZdDKTrf0hNnO/VVK5ohwG+WpnNDyZVV
kLXzoMk8bhbOKfRRCKx17JO/PdVi/ryXmjY2RQv8IaSL49eROZt9udJnprErZrV6AQ9byTKtctvw
PEE7F8hcUDb/Ed0Ez7AbJWS5SAFNMXwuIhsNNyXt3Kc95bZ7sFmUvBraJ+kI6+l/HIX+Y5gfE7Am
cgO1OQsdwH0bN8hLITspVz+99DsVqwqDreoH2othWPpW39NYCffRV3WcDwA3a8r2vMuQnmyWVLBZ
OJEtPQh71//WnwvHxGljE/rC7qDul1SFme6jjien3nTUBpNc7fMNNjqpPPHEgIiHEhP/qNH3U+zg
bmQsg+eTIIL7l5aM0ZxWmS4YWkbPuG+bvERc271dzoPDiLJsCS1neH1ty60B8Rs41f9XuIc0J8C0
W/kUabNlnsA8JQPiquyQ/bdP54PAGnB0YZhlBAsjyOpMGKlub4bXp1WvYtjbvQKGQE7KiPigAiLA
bU2JHsoohpS5RB6UtOXouI9mJ+ObmvmNMrAizwFid1cSMEfQb+nnmifq26hy1MC8tStbcwmeGgz/
OMUqWITCpF8MMuYR/doV48VNi8Z4cqEcmKIChVrcmLMF7ygOBVd+7h5TSpcy3QTSdN3dANUTqp6E
UER0ZPaYANqcp/sDARNm9V7xOoG47MENb4zbutx+iwJhIGD/4sLDb36YG+ru0tUFVqPssmQBBq3P
U3QNbBu4qXcGyiaRj5uTRFLLugbxJIiBcUn1tUIQcOu2W+hhWW0BDy3HdmsaMMP0+KCYG97nphv0
tU3bu6nTVOFntgJkYk7Xb/ZG5jbyYbPKKpL4mHvmYRCEm2bRM8ecRaspmZoh60ag9IiiB8k3L0mG
KQXz7tjHQ2Tb8Xncz7aFlY85wVtN5gHYQJr/SL7ytFhlzBc0iF/TizNgGxcogezW4Fc3mRIFdzKH
NtCSWO5Sq/5VLxZ5u716+x+gGQ+pGYQuyys3ss81nwS0JQLiNhlhtpIJdhoaE03ckzzUoqkawy8m
7QPwzn8Gwe3gFAXAu/TiNXNnOLod5n3jQLi5iixXMXwYcNsSx7G95ADAN8wZrqpHRHFJS9YGGpZc
raHGBi0yRx7Ke0v1lsyZ9oh8gawjyfDQWc/teVPpow/fjwLt4sFVm1MApH4spx04WPIzP0haE7UN
5RgL+nLJBxxc2UvdrOFEG/x/6UHpcoPL3pslks4EedBk7C/bHPF+IlZOKFjoCLalr5n9kcAhT78a
B0eW5xZ8YMQIyOwQfN8otCm2mC1dlKWtOGV6QDcLP3/FIRnRZIO6fPn7uuHJ9MQ/bnNWjSSk4XrR
sFwoH6ARpXoCi9PYZ5geLw2ButbYLwwsRDxOb1hGkGDEx1Qw3Yghk7c/0EAcOxnnoJan3d78jgnR
RkaXCDeFdaUXctwNY7qjTk3OzqUcrRzSa9QBLX/fK64bz03OCLB6KS1Kmpp+V0hI4sJ39OW+lBPP
4BkrRI7q5vJJ6MkVYKsddjgriF6Cxg5h0GcZmZ8lgP6ozo1V01FyoUYj5Uxt6RHUTg1vcGyJ6TtI
Ta+1O/Vy2atYhGqmvUbGeF3PIlhSxux4X9t/GnW1ZjW+6EJO6j1xtV5U9NpTqWJyqthKywcAXWCk
/5c1JPxx4APTcDx8Tvg/Lm5LlWc2R+1w4R6ZVwY/qUMmG2PprwtN0Z5iT/x5RAt36K+ehawWMtY/
yAl8suzZiiLUzZ1m07zF0P+cd0M47yRUfnh19lirLX8Z6UoU+o//DxpsnquVrHEU+/QegqB9AHFp
cGOOuhbht903IAe5O9DPd/X9uRH2bb7ctUzzYlzORt5MTXEWaB1jsKGaVKA0ncutkaN8MSphtGQy
WaykwuvJVDli7WnKBMkl1f6+EW0i4HqH4I6YM1/3WC4BleXgN5elyPzTeznM4hZSgCU9dmtNuKAD
VEkleTBfHEuPaLawAZmJLKhFbVO7Esw5cQs6rpsl80hG92+xkjEawQVEmKdH31CqJB5jaP/4gAJl
Hep6bPPxCnjlp2NdMvzpAgEWLok4oU1NudH30P5O85BLoqAMzJx05f6Y27H3nAX5nvTYXH+uUlF4
jFBMoSAS49GjzfnzkHYc3+s0YsRTgylInw2rjZwBgETwpNkcqmvkChDhAfOTspP5tOylOAQOTi55
x7NIX+wnTUqesLtpIUzSGIBFDV53Rbzvf86cAor+kgiwAAWoee96cfpp+MLPT08gENoCgxPAwQPr
YfdbyPkEG5NNbcFKFv8VjqhxadqePo4ejRe7preEjeZX35TTWc7DCyT7qfr6c3bSNC+l8pXUHA4T
7ZJesmOT5TNkhx7nWdbj1gWQTzgZnlV0D3on5c1qAhBf4WUWk7TKZv/IR9JPvTcP+BwNRx9lCf8f
TT4bOgcvTNAsuD7ihfdH9glPqjsSOWJ/IW08oTkj9YeLU9pSpBMkxq5MQ4Hj+KCbFq/4LMdFvt7q
G8sPPUIl1LFdvBmg/j+mKZrSl+xa7pB4G46PzTdDnEnWfU1K/21My2kQmXZWfAy+eihlhOb66BPq
ytWwcwZRtHJj4FjsryE9UZhBrD5nO6h9HLziNg4P9fPXCrvNIR55pg/YmahSm6NksFR4OV8uGgo8
j5Qjh69ZSrjdI33ZK4GMY1buvg9tZiIrH6wj1v8c5rEySMGsibcy+xHGT07XiHzX3tBnXp+10Is0
Sl9jYKCfhC/DWFnzSCd/sCMhu6AujfGd1dUUjGink/ELhyEl2ctp+Pv8/AVF7oUX0NUFIQTSj6Oe
S/KRoHmFlHP0XfB9sfCjl0rfr7u+cIYoOxIKvCF/ETYxKeK1k91P/nQqOh4ZwdC9KtN052hj2AYO
r+PfmLVDqYH9K6joE8oOBI1lx5Ks4HbtvFzS3l7SiUownhhEVCnI+wCHrX9e1vTaeQ9E1Ob92KPN
wDYwfM5vRq4/zYFm0POIfRk/P+5oKltNlAeLtOjDpAdjW8zzNWJLzrU7iWkjfhUR9XfcgTIbWwvU
Fr9Ak8BVEPuBisdjDZER9Og5askfOl3/5sThlxOLv9ASlrhAWKpTAfHGCAsXsVNYM93htMvqK888
FJgNrG3v08Iae6nEYgV2oUC/2ICCbJ8bfzE1deqgwx05T16PEQncU7zapPc2p9KcF0NYcW1356tq
SiRhaDksXVtIFR2cWTWSJVXQxySMJ/KzIUo/z99MEDzvemnRTrOfEmTP4/0PLAqqxoDxjboBZOlE
80HsY7Yh0ovl4ijcFEN+i1Z0gMSIaOLePD8gUJVmvWi7WfdJKHTf9W95uTBDmYVw7N9HBlbfAkGa
9ME4epIhRlsj8xVrbP3/1HDRw9nZDXLv8k2UosQZjH6beXWuY9JuziMiukPEjDWqVcBbUoLbf1tq
Z/hfeTYq7H3ELpj9vwnAsAaxMsW1DD5JjQTS1d2E40xxkD5hSoOceFlRyKNEmbGULlYOfwk4N3Af
vubdfAgZtGtVnxVai50k2pSxnac6U/mp7mwRTknWXTc+vN+rBDSwSzWdNww0gYfQ8WVGbE7lRiQ6
QFAv+3cE6pC3jcn3JKgUJHgoa5+X/vAY5fXCmodISaaGrqGam4xcb8xn0mBZk9Lqhaf08sl7NAuf
brk0wgcg2E9r99nVVXnUGhOxkng/SDc14E2U3CKlJ3JgpaQX5nagUvao63oGOVbCpioRoTjFTHNm
XcbZ/GmTfzEYik1vHxXUqhlDq9VGzr3OWI+QZVh7UIs2fGtfhB6HL+XGqdDsD+KQ4clc7lkS9rVu
ALV3XkEPpPYrh21xqRg1c7MaIdzCrRxXun0wGgM9ob85hDlshfVJ1ngu7DOPPB9fBg3c69SHUl/+
PwR2Ol9E+id/cVRTW2NZntVmWL/C7WBn5CK8HMgjXv13BoLYjtxmulP3io54MMCP5skzaLMpCqNr
ILmJ23jLHfLqVWGs9qTfShxwwS05W+uIETw9TsTwgwbnhbUfye0z/qxjr2/sHiZf/8NwLFi5KOBn
tz1o1qg36kvZHKZMGngE4ySuSJl9TLnYh1hIDFkZagAcp0+L3RyaINfBINQ3MXXPNfVo9ydwETW5
Hw2iwFDC+NYF8jRDo8iry0o8BTwFByIkDDw+SDazZbxDQxC/8GRcZICzsTOEDNDczRcTTSxhEBqj
GyJcI/eFSsju4HCEZVL/Wz9plwkZLZawSV3n16FOAjan+cxrXVbXe/8+hSn6igJEhhUYzB2a6ad2
IotCvvJ5V4cVnUkEaWx0qypTn5QN89/hXVmHH8SCaYXP6+yj4qq0nSDj428NPlYlJbbujeexNMCX
3zZCZZw2DU5x3I/xU1gVxStvXTFEAwa7K6AiMRuLb4R1M4MsgqBsrjk8sjnms4rA+r+LSafUVgyP
j9/W/R3F3MrQ1o/IxruZJmT22R7JDXzTPThPjlp4/gKHH8KyP/fBMlCbjOi/ID2eqz7w0TR8WPWB
8zbj3o1T+b2ufkPqVXpIPCS3Wz6IKRnvbnIQjEL4Qr8WYv8gry1uEkiSMeAoUOgMPV6zOD8ad4/E
QCS+7jvI4EdYYAPBZjWOAe9SoLzsj4mQot9OSzPq0RVHn4aGo+nYYL/rIAa0+dZGV8jUxLwSneij
FncOh5CfN8bjYc5DgnS6bOY9O9zQED6zGbexwCKoUOS//t/lMWfvsvzwzZ/3vt0P3bxoF15u4/A7
KgUQFXZmA7y7lkkff7qzAsPAm1UGZOsBOuVRDXavtoRcHfbQVEV9zBzST4f2optCfGR8u0NooL2g
6uJnSN7b3hcGeXRCnYz6TR7GPw9KHqS1GfnJTQbjuvi5WnkktcFu5I/jdAZEUaf0caP90Wo57QVN
GP970JLcs90NN+ih9jtE0rzGneT7fFHx+6Pp0RE6n8kMKnZI4u0YxqxJYs/LNhGlQP/51t9nsjL0
cv1D6y/6WE03DT9z2vUmuWls4e0TT5+GCGCP0leJ6a7BchtbVkKZ9bkTcsSY8Aa1UuT/XiOoALJ1
8RXTMMP4fm0igDSy3Q8j97PqfFsc3CvY5EXPWcHsrtc3qV22Mqb7G7ic+B3rdRpO6raH0+rBuwL3
k1UBBl8zZ0+mQ+L35IkJ2tXYQOdeXSsgsPyZ9uwtKX614LyohU8p1RQipkK5Hl6c2Mn3Ck6vQnNT
zvzTP+ouh845HFe+7dtV4ibF51XdrynjGVZX+OMj/WfqMmOlbeVkePZcQ0FRHfqlU5ibI6Jmm+z4
LwKH2JhfZAYqDtnK4kSHbnrrQbdm9l3eeeze6B/39g2UnLvcp6pNqMwN/sQQVXOen6hnZFula/QE
5ParoxhbyfKDE9N/X3asaAZaktIXNLDMp+T0aLRyPVrRvTftmazxaVzrRdO66vfYdXeFFE54SB3X
nOJz+Fhc+nW3L3fdt4uVU5R9IGlmnU5lRNclKB8LBMstNL5t2kNKAIQFb3FWHcP9ysddSw2N4sv7
xPuB690X5pVAHZwqYJ2MkDSiP0o+WQZpslQyDYaFLvYn5HjcvDOSiTBmUutRXrIzKdUZHAtt58D4
9xmJocbMaVdbZwtnJFX3QF0jn2FKvl/FumkpAwIyI0BpGcCS3oyQCXRpOw3ZuNNPt/nEkx2CYwke
qg63r68ADGJIhF5YJ1m1A9OA0J1xUhfTPH9ucgajvlThIUfNEVyjXPs1inAsv7Pn0ILROlF79ioO
5OJax2ehZ1lETpL2advnEWCj/BnE1K/HlNFwCjrLMPtytZn1TvDtCg2BOhsQcFCGQrf9dFPjVsCl
ARTADPDGvnLstvhjw5WAyiO5s9ipjaWKFSorANo4y34tspJtGpHS435T9cbXNXbdHm02ybvlgKfE
EURHRPRHMtG6VV6tyMCYkcfFfpW3K7bU7/yZRkPQPmgQO+IqbAZ3j/ZaGZvM6Im2orI9koZuGjQD
0H40pN6pjZ+NcSJbGuir5LIaQ2mRBskEI+pUGmVEWnrzWBF6FaK8ll+YhVS3IdGJ9PfbLVPG5GGH
X9yIni9U+EL1KxdAISSd4grBAn9qRfZaxJZEpSie9pRXjpGU5hTX7QvyFVd0s0PIMrQZwYzx/cE7
uM4wPRdJyUJnRIWbPILxt+oecgUSK+VB83lRENA2TuiKYKJ7kLVwB6ts8sgGLvrp55a78U1+KpNi
OaD6MheMyNwd/YwyiLwM8el9vcSoN97CzpjDFNqZPIoED3CZG5FjxVPiTYXznbMBwkBQrfuFR+K/
qdhbOlG/09ycezMm/hXGECRMuJI8ebAW6FK3iRh+133awmsQcJMpIl+2pvD8/a9pi5/46VdfPqeh
RXTjkn0pu8ywfOoytVusyhpn+zDt2jhGnsvUTt00/1WcnjTTVuYuc8R+MsL0QXG2EMAg/IZNQt7T
v0dSuFaZMYu/8U6zEEMM/hy9etT5T7nh8VQmYRDpBerxsi6TZ1hJZ7tkATomKIlZP8UeZl/mhwNf
H/tVG9UXCoRJ/cR3lUqA605cM5CngXDh9hgJBMmMgVfc5Zv1kgvxSmOGI+tFgrTeCWYheS06+cbJ
y2Ig/CvUzV2I+yC2i68J3QyPrBni5mbmtevBU9o/Bx9Hrl+fqtzqzN8g5ysiN52jZckIBmC8xtpr
aD8FeW26yz1C+tUdYQoBGwYfedbDCE4UFko8itclxqRiHlhN1OhtzVCaGusa13q0iwA5ekFK9F3E
SH5YNYw7B5nU7yRQSu9vsgUbQDSrP54utWLNgUC4K4KX3HL8A9JDt0HswWdun/s60fhcUYd6bqxJ
rULXP9JqSzKjAA7r1lNVYJYQEoDFjMor8nq7z0Qg5wN0QQZOoOjXpTcL4QJMAhusEgWdBcYrxHNu
eBTeOHQeaFbd9+4tBLzxFDwefMOCYviMqG1z/Q6D0h1+Hj5RBvw2QIbK/9tQ8+0AD/zLnB4tAoCL
LeOZPqAUVsPOKgUcQ6Sp1xwsa+YbxrSBWKgUPS9DfA0+PcrAsQdsUVO5QsBQcHLq6lMUDnZSiq7Y
grYRO+hH5vCgNCtuQP+Skxk964DjDisB35THLYOSsD5NkRCEMrjKTFLsAQF9RehT5Q42ipF7zi5z
QKbaQDTqhgyxoGuAYo99qxPmhbFgLEi/Y2LDdjEubKGwDT+dZeiypFi1/mrq0r+SO8yncolQPMIb
mm1twLxR/rcquLRheOsuOtkLG40v9/lppAm8Jh8t9DqfAUi95w1hJF1CUZR0e83eTyMGKfhjuSqG
WCFT4T+c0vzq+0yhBCGENvtJ0sCRDPACsOaiqApRUKTB5yZ9emfhZrnWAKol/YikW3XadssM1NoX
8jhD10LXA0ermoVl/UJSHnlq0BWgEp11bgJwy4vHC8P4ISneL9nCH47JLMzWzVDDNZgALIOPOWpx
jr7wTgWuLEnR3REC/KIQFTIQ7KoN8ZLAPGBhqsg6Ap2huYjKhVum5TWZ3LBEATaQpiMmM93L+pe2
G37Wmu1Ij+jQYjoLV8xfwhOztW/e4b1E9Xu44v6oDtRxG/tkkXfO6lSCOohNsE3nVknyk2dEOd5y
a0zZo0uB+XwK/TiuifPXQxttt9Pz1W8ds/FynBb/MeZ9z6wiFqa1dU9AOwJgWsPfZNvak9OR4PRM
P9I8xhytV1C2SxTnVLxW17VUZ6eO0pWAFIISJcazuWafgqMWPKj2M3AQUUDynmaMLT5DGTLs28fU
YRjBVjDW0QrjaZ01L5udPckVgrMMMfAajuH/UyleZYKqize1Rf2rtYQQxst5QLbGIz+b383qTzsj
Mwpr7+r+yKlckgybhsaXIWdb3GGZWHM4AUDLU3XcMojoR3WMZcOeiy5948U/Ddvl6cG4ThlPk4CZ
8DTs3plEaCCy36WzaBtms7staBnEdCHA+q9BuNWuWGr8yKQT3BuvyGoN5leJhaTxq+vQ+c21zcOd
Fc6u8zs+iswEeeA0koNnt/j9VSYVI4qOO1EnQ/o9iNRD3xadH4oJAo9OfqTDAojlArLJMlKJd0YV
Lxo+JUpq88yoAEAryarlFxkB94hI/arQkbw/WXFEz3OfwOe+psNFfzH0S4biBapx8xgX4pyYqyIO
xsZNYjsbHBLU43QAoXxklnS0R+kbwb0uRhw77/RchoMi7WDiQ+Ngx5wQyrjfDm65X8UiVgEVPDAh
zHaucQNd1HZQdi2N9Nm8rcgaKh/gYx0V7b+8PCXCC0zj0tMeZttwnjWFV8z4PX+LGK9ylsFlgYvy
v73ilfDUGokXhep/O+Ng6QY7vicHpFL9vOHmOPJtlFCo3qE2A3UYzeYmiG6X53no5964rUQ1jx1t
VU/f9kzT2JDUsxEJYkDHwIwhJiOQNDOE5QtVVgTiLLY8rugXtaNrhEinopUTzUVBd/utTkxfICDA
SothN+g+icOcwYSb5Y6h8Vp4kVaZvCSe75k4Y5lCSsAxUjwd0qMlKkxu3Ro1Ltp8dle2Aoe3/zRq
f98r1urQo7YbDeGH36KSe/On3ZkXhs4mRdvpQfsxKWeD974HpfTVtpckg4tkhbAGu9fB0E5oRt9J
LUDZGNxgWctnScLeQXrokXDQkguPJSS38EvzRDd5Fo7FO+gkZcurKFDyJ4ZOL5Xy6JlABEHdUh92
BZuqgmIQdLiiHO+Eg7AskpQ5QcnWNXQ25QJ7qLzHe0Y8TXLhwXXMpltkMsnpQcjlRGZ6qg2z+Gqu
qSPcVY8Qdmcan8kw5ZNuDhpO5mDqMbsjfeRkY19v7cgQDRukOfysRiClq29AgckvG/ngHQvG3eh8
5ou00NCQ6N5Xp9ODggIbpoyU+mrF450kZ8AQISfjfBRuV5MMxuI+eU49XYXU8CFtctXzLgxacyrj
obTWenQq+eD67JJSW//aZTNd6pW9aaO9VJZ0yp/lSHeSv/xYRd7Sf2xP5m40s37YA9pyTKjkNAZn
LXwEQ6G2kQjwrsRgIXshh55+W2iARrOZC/E2pE5GRA3cPhvxojE+2jUCl+5ImT/k1QA3tBZq63Gz
vk9hCKhyc9XORjw0s9B+Ffk5nHhXW4bV5/Dqa3Y+TT/H6VvgMLFy0qPRu+3hXy0rxAmxgcJcC2Z2
5lqnxGvA6mGRp09xHyrqswyDRpjSlfdwm6Z14YF1pb4uRyoTLVPu4tj/xf1NGsr+Yr7R9tTMVFlo
d/VyOm+D7f1UmtX+AB3ZxXsAK64YtjuCPbz0Utjrvv5bVv59RtWsqgBa6RPjTXwgO/0ybTWFt5yw
wsR2FPKASQhpntbP7khFu1+Xe97YN1GRSf0Not93+kVX1wEWDGhbfeOCLXO9ALQgVu0vbr7UbbGO
MhVUQvC6tgySaKybPwEG8vuQyDYVVQiNnkYaMwRN/V6zkrTxcNeVKmTLrBPKSs8ZHsitv2yUn6PN
DbH0foflgAl47JuXhiCaFF/L5fMWD0trmG25Mg3bRJwDu5bkQ9nR8OR4XMrRCWNaXymNnjWBlluG
AK6u4obxLINiogMCCmTAmizRkcMsBdGcAnhvdzQY/BPIQR/d9H+MO9xsx+/x1t0dmjt3diHW9/k8
QYxTP9U1rqrG+45fw/r7xQwqOhlvyN98P56h2u8R6v+XywlmWcToH4l/Y0xOob81EeEtjy5Hl+gb
wLuBqfUgEiR11CWc0J9Ac18dnOegaL//oZAx8EIzmIGNh3Ad6jeFLlbt71vW8q1O1tJVkyLuxz4H
hS9xNPb6Aae04KBGFBxcL4KfvzUPVq6z5NM1jIFwx9tFG/BrO2jHUzxYtEE5+GauC8p9L1eE8N2b
kU8d60bHcgRbIKFDHBBzbJv1aJ4DSNIIfuo7AxigdRWKtGMRcNFtVYVmS2CHwzIl4PGnJwxoKtfO
7xqAljZhwp2FkjsmaTwioWNwm8Udx7V376Prn5OjFzOqitm3BTgVGwbGjXta2TDIa9ifWo1l/+I0
++/rsdR054KWIQy4n65Rvja3tKEOkFAJbRF6KbAd54K93sHOgVMeFCglqGoER8N8Xer9C0Q1BfwD
D9GUvFk7g2ujn3KhyvlWNy9Y5plY32LYvDwwQiNhDuw8yOOaLcV95w5nX7SXfC/YLJrHtplFkWyU
bE1Bk87Ne1bpT+EWEMSBzjjfZ+H/ciSFG8oVvXx+PSeDDOGGsUZFqDfEOai13YzGoDkbVGbdWOPh
PLa3yUwPMi5VvcD3BNCafc6O32uBLgr9p8mV7btHCjLTcuk+ViJuuBmmMHmqWLij0KUUzD/JeWO+
GvsxfsPqP2iF4pXZIczgCHBSPSN/UmLUn/znQ/bKsCvXz1fJQ8zTHL1FnuaHLiffG6gIty2uzWzF
dSgFrNxGjncHeeAgMC1Z+mv3Mu54CEAV40gJz67uziluKn74RRLz4QB1qrPry+200erZNot/+0D+
THV6eKTZjpRr2sSaLtUDshE2wTeg+k0HNCEHXZjhngAR6QFZzGZzG9962E0sJJCs8qY+XDJDwNow
i+ZujZQxSS0qDYAJ66SFi4+vYHMY0iKVGgjjYpGDDqR9loDomiLFjk6vdrFs4s51KsqgHCZzv6VO
9r756N3+fe3JuxdxR04+mBVSt+6dsYaj9MMz7c/K1Hx5TNcOtpAvmW01dCjo1UGDHFRsj3/Gd1Iy
AsDOUZdORxuUArl+SQUgv8EbFz/s6UZK7i8Fi02TSpkHoXrVx4gsK5KwpNTwQkMikOkEyJ82y3a7
Hxk108cuNRxH5xUrvNolL7JuSVR+pWWOsJWq8aY6EZzMZKcnqgMOQJrK0de7KJZ2VY5qYuac/g45
+m33tmpcRgcNOrFPbbS/P3l6eukZNBpFa3E+xNNDcVDwe7sTo/AkUaAlJmM7t4HXUFlY/Fsn5mZy
Q1S9m9fpf78aW5Uw6cRSZ+Wpq0kSq8toXgRupi3WsuduBUGAqJUhPmElUk7tNyC9hGcbFer27lJg
y8U2kmDK2AQMbk2prGFMTglYO0LNwzLXaU4SQu05DgibJ92cexqR+OhK4H4b5PuiX0GiV6P4Q8Fd
3k+AJKpX+n6yQfZLZ0uClrCQmqs8JCBEzGitvBjEBojmwVUbDcNT3kaXfUdHU51KI2mCtYvoEraY
9YSVTa+Gn71d6xvhBVyLmFMe7fZghN32VlMhEgg1U1Ue4RCaQhR784zg+/O/v16gRBMAEi+hifZl
c7SeX9Dp0qxfEkhWa+ssYaG0MYdOLsl67CAUwYaV/6hwDb3eIfn76NVC8VCA891CnozNLS2hw446
jXc5g3ZFaXHtamRKR6B4ez7VpopNIovM5CC9cOLC7/+MY4OiRgEggKdxGdszQvAVbgK4TyAX+KD5
2CPsnwgN3+pQ1BNlEOZ3Xi5OY64YcTegcdTHdxLnEdCcj6J9seQfVidCpLhWIRFVKJw4a4mOoNfq
mBEPQjCbDDpMMgEIDg4aU2kpfjrc920W3O1GrhDKylwpshotb3yxNVFRTNCkCOWwmuvJa0oxVSw6
wdxtUwsrZiRnPbqOENCl8zJnzB0QCYBqEglqZlGwi2UkYmTfu3HuE6UPX8+xIWVkt7cAmoBQJI74
ByXVW8WNw/XbdSkQm1iFutQU7rRDC3w50swjbH/GVVv+EBLh5aBaA08QWgX5hsZwiW0/4eKz68r/
2HA1S1eStzAtAiFPCARoc1Lafsh6PnRkP8J6y0gi+gZoKkxlHj02byy/RBKb3SK87dZDNUctE8DD
WNKUVC7Acs/xmbx7o7Vg2bP0C9i5mtrwaukNd+MCWM6IyabGhR+LbuitVzLYYvlMmc7ZpmdBSDOj
bwIfrOGK4SgVQbMJmTCe1cBo/9CMK9hfo0swTAMbDuf+23ia1IsM7SsNlPJQaS1IRa5WyimduL1e
RFEpS/lnZa0W6rUyXA5jC9rrogicm+p0WP8cFrCO1sInfXS5i7fFVlKRfIBF2DTQLpljhj4XbG4Z
PAYUzqK4KS+DRmOHmFdMbWZ7GP/uSNcXGSMwUZGI7dDvN7UD2mJsiAurLTyiRYCduXPJQUuymtZb
1JWfWsa4k7VoDG2fM/nTHakQC7ylicMQvppvvix18Z6CUpiHuV4Z7zFJtqWdiDg+aSKx3fEAjw1Y
xBypuyO2Ynp3PgrGOeMRsA0m49Zmw0tOqXOMa8xSgqODS8kVxzesWUN3+4/iguXBqYysBUoPXZFn
s1d1w+nWze8TROtRoQ/PugRUy3g9BURIGnF83YtoDFTABHo8Cqe4tTJT/9YbbqA+WImH2PraD+7V
a9j1zZDG0ixejQU38D52oBMO66E+2KM1aglpgYEAu7P2yNJgmjz77ev6rmn51jucJzsLghGpq6C9
75J8NYQzMJqP1ovLAAaVFXLYBF11mftK0NL6Vna9jv3YnyUbb1EgMR8iS5qnll968ZyskUZnfIjx
KAre2Ku6m5S9dp2BsQy1z4VWTw1MpMn9DUNG8sPz9wkxJSM9xNCqXfZone6zk/YSqxeUESsNiJXz
uMngxPCsRJ10lOCOLZp+W4QU4HBNqEJr5g/Wj64wanB2hLU1RCcZBYv18FWn58tFnER0CtVTEPfV
cffS4LNva4HtGAemjyGy9NerWXevZh9yRJHNfzrwiBjseYyWpgoLNEt+GmyEM63Qqc/GgT0fsOU2
PfRN2UzjYT751jgrZ53sME86ptsDSDVdT2LZ4/wlq3uQwtODj6CMhuXX5YkTORlPFoC5M9+fqu+h
ciSQ8jt/fC/H9e0GX84qCdK+HjOiOV0bhTS4HNYL7TeAbKeDKF3h7w4Zt893wxOCgozFRCfPQohT
CPEkhanOrQFx0++dD9W9DW6hHKwU+TTOmCUaUmU4rV+ib3sjY5zCh/CIkZH7pliwmKuNMkapMo9J
EIJKNGtLaDbQJNRrbSTaJ5HwkCu1NpNeaeclefKUQ8N0h1Bs33AgHJKw51z4WUHxtFG6+F2bn5YP
wgxrBWygKGxjrq1xof9JoYVhf6LAsrS7D7p0unQ+qBqew9D27izRK/slofDbIIZwatcvpUnVqJmz
IlDqW8Vn6jFxkvo2vdzh+pgd6iM+BRIEkn6OhABi5ayQd5wGj9VF7CSQ/wXyaWd2KuW6pBFG/B/x
zUNHqeAGujgliqE/CYgrIeQW2mtNbiKsro+fOvocVNo605um2HFIDX1gE9vCOiwjunL+wJYXJgX4
Gg+UHO33+VKu8PNk8CBjRhubqNrF8EEwWILzeDMVlzcy6O5yWqEylDYKgYU5cgsOy4bcmv5PLVH7
QjmaP4LK+VzNH96Js6cYEpePN1u3AzOlAJbuVNYECC1SrQaXY2HJ8/3urGtfM1pq7XGG9DlMkulo
F199ns5uJabQ8GLdHxw/i40xZ2oEZYlC0xDapoYnI32XXd+gHorvVX60t9seLPjbQILSeSN6xMJ0
y9eIKRrWl39htWT1LtRH5lesVHlDlKEmFiIqhR4lIyxjavpi4zSf974NKEIOy9zGflrMjcHeGyiE
C7KrXvyZZqyNidiccEeJD9/E27fra7Sioig++MQzXYP9//j0p9WVWQJCUJe+fqkVwipEtLacOw2E
6/jy/u+2DUoqqfWKVM/nlne3e+CQG4braVrgx0bC2cQKOU3YsEOtI68GmWGa/qH66neK8Tn7UKvQ
SKhTmNtiHb6UDDW3aMJXJOCYo/HCox6UMpB7MpsWK/yx7zFNJjy/pD6PuzMAZS1inePHCVF2zpfE
ESyixQjuCJ00f5+GhQ8TZTCuYZapb+3CWm3SQnWlCBdh6SxhSAmsVxKSYJ25QsnMXLtQsTCatIDu
KiWdMCCVteA4mpt62J1TJ1feU73BY1D99hwmOHvgpw09g8+DAR5cWYIRaqdTdt9vIzbpmqbdoQ60
RyFiq+BBplRWbx1tB+TGjnzKDJXzuc0pC/6EeHE2XQsa3z46BphLhcAq+2ekpc+BzU7SSU1Wp3y6
z56oVfuH2z3i5UZKK1lUiwJFJDhJH1jjSfMCkf0bqlRnkE0Tw2+boOaSVNfhiGkUqIjeeJgzRI9s
sjdSkkqPPKa3jxCigsr2Yb6h1D22+/WV5QEdLFYCgoDxePyu8I34kkXh+MsclRwoz1cMJ2C37xxb
UNhkwsm8j3BWAbvoXOdioSyq8pS+8runJeF4gBZG7T7Vew0GDt8/HQGqFeWQ26wtl3ZaD9Jm8IH7
Pc608Op3pzJuSwAi4kglxQESggaqxOwng0vCTI7UHntPDO8T4ItthDpzB0JFvBd3MGV6HwXL+aJg
+8/SI1+takqL5iiv4n0ZSMP+xWiY6frjM+b9ILLLL5mqTv9IWmNb6izP1Imn3ePlSx9xd7prba0T
g5d+i1bsBbQ1u6WA1+CoEe1XcUhQJjtz8at+177ngbIVB5KZ4D/wmmZZUFpKC4O/dxytvXX9h55O
QlduNtLWFd2gIxO2u6SVImhwYYmCIXL5T279XojqbkCaUPmqCdI669I8vbJjXdkbF0M7jTTuzbQh
kvU2jVaIPfcIF3qMG7m2nphIm//IOKM52FX6ltHsVkAn6mjgSa8zyxFn2tHEGxxGJToiKz2c2h7g
B3iBBqpTID7YY40qLextYQRHZqpQ1RAB7ecNS8xwTMXFozc5pf7nNu17KO86d4BwbsCffoIHv6i/
m5ckk/oN4MXW4YtnkCgoIqveotOXsgCxPZQ+/6OkHwk28qxR+1Hckxp5EGmVsdQFChauJIok2EKj
pzj0UcTdghvOjmB0Wo+Ff/wvYGMaD4D3jilCoiTHcAnUDXGeBldYfE/p/Dwd4CDtS4NP9Kx8CyJz
dL6dYCB6now6my/Bc+j/PYw9UjZUgv+KzmFj3ycpvGJhfZgxhICYlrXiHDGte3yBgUsZLgt8YrWo
S7D/p8zFWLqKtjFh0D+ju8SBWOsRTGp9jb1RmMfY0i1doUJ9syFn1NgazS3MY8dhJpf2YmNQyEr0
vCnvXVOzO/+3FTQoM2ezJCsfr8O3cF3Gh8+g+km40lZLdMP8rBS8ONc5FLCWFnJMGEroM+SlBIpq
dlGuluaotTcMKOuAQQ+0dPQbzTSXgsnfz+jXhpnEZOweAsaaf5qM0UT6mgKTyO9BaxTEkqL4o9Bc
NaeoKuOHwgXNay079hZF4v9fs6r+GtRYOlUIyxGVoDPbtldOQg3urwn/iPPxOSPeOg+zgEOqlwAJ
4KyjnFRpwRYVFVWZ0pg6ujwO4ETTt+60+qw3+wMtQjs2upP2h7roSEpH87q35q4i01GZiVXl/bwO
VQUDNuBsQ61P8zxFkCQqUW4TfjH2LRCo6AE8tMN/m5qz00CEnYbOUs1H7ZNoRX/TNyqm6Ldb9HtX
tAGm9Xux1mEp9w370HCTUIoctCCGLJfCu+csg6PY9s59e7+/yUDCwD86KXYI8cbu52ADaoMR2+Pa
knBcQ8CbQIReAgt8nbIJBuM9p+qLSXJUuJyxbNqpXXFPdqYDdkNQF6s0IllCw+dKdHreZ3wjVFoj
+wgrZ01VWvSbA/HuEhUN6ickwLvAqP3EPTCxY1uYyE6so7gOMLo/S2DLjkvOyp9UrDEoh1x08fvV
tjAXWxwxsyzDR2/oMOPYoanqw7kryDHszSI5D9Hx2fCJAhhvsIiKvxQmSSP7p6W1uK1oO6Zefh/N
G2XeOgx5woDRC/84TNrYOcbaIMUNxr3lZUhhhDLh46g84bANjfznRGeikB/dBeEidVjfg+MkPDIL
fvUF8KFM+qzbF5qDI7GClzTjBou7WO64/W1P/O92HwvpBCAb3O9Z6O4A7IxurNO/AmbzkCxwBrdY
fKC/MZxWbJNHjCLW08Vnd6+vJvvthxbVSBKfCYhE5zvZAigXLR295Ab9H0NqpCq295p9vgLxXFGI
ZY1QB1WUfit/ngOiyNgzeZL6Aq/37H6qhwybXgPSkR385vnlN7UkSVUURoMeX8i4o7kquFVJWTQl
Ey6mk4MEqTL2RpUX5XVx5GykH7TfIN1WrpJEM3Ugdvc2wM1C19A2CQsZ12rKlmwhzY8RLpY8SMWm
VfE/eMlGg8oVCASa0a7t0KowhkMgzjxOLuAoKjhCmLm2RV0/vQauujBJt0+ryP1IorRvCMR9U8WU
jiO11BtT/yoGm/HUYlCRnCkGwQFru/9+F9iVsLbM1qCBPOeuApNvj7/g9roE1qIV0tiOCcpvhkek
x0q2ry44aAIl+9QN2lSRB9aEx79uZypkOxqvgFM8qX45PF9psTU0Z2egq/gUDUD/51kww+h0+/dz
uKA2+M79byAhuIECTid8VddYpQniHz23OhV3RhULLccJSKqYKgZkqu0ruuf+x+GAovVIHwXG17Mq
t6f07scwhE4N3p7EvQWzHYeRkSyfmZ9vP+EwUaVh+dfg+qvzqc79H7RWj2ewHEK34YeWZRt+XUNq
r4FOsg+oJ7D+tBDw62adq/h/O13xQ4IndoQmssMelrr+Ga2PEe48NbAIWqPyWixSC4PubINvuG8S
Mube0U/ikRel0mZf/wNOQM5N7wI4dW3PtfulpULxwCMlN/aSRx+tdFK6U+sn8WnDZZtyIaaCJ/Gm
Ag+Im7R9Kd748OTvAK4MppJxeU2nN5guNSsFjx5EthhLsQR/iSk61SBCz5qiXY5XfMDQONzxa2vd
80xJP+2rqEfoJyLvy2NzF3XzUh3afGNmNSmYYHBaYPQw0KidovRtKdtMQ0rxp5/RnB3HCPuF+Ghs
qyoVvKeCIRV+mZckEtRX1e1ShKUmDI65jScdD2/qpjZopahEIOzFmCmPk8cPKxLgqvBFlqNK0IYa
/QcLwrhXVGdkb4iAtYH7PO4ePNYCkc8hjsFojAiYRpa6AHgFF1UEa24QXZ+4euTVzt75cT/Gou9S
QI2BlQD+LC7g62t8en91l1qPl5I8g6jG/ZACFeFVqSLJUYj4PKvSI9Yiwch8xJIsefdOXg9DziI5
qn1rlABzb+xWFRhRx1vbREx14zqJ6wzK/64cltKENLqgZJ5SG10HFqSkq2dExx2VfcFBvIbCZDZL
gT32CSdOAcZXCu9xyUkbTR6nUWj7jY+YSgNqtjNnLHE2j0tY1XXnTwG6qQtcBGJeev7zro6NK1LC
qky9uggiLW2Qyn0Kz0ueToHtFJFggdvq01CgYTcMfqMBu76hmKNKrh+Ow5N+hRopFO+0QNIsr8Li
dk9/cDKt1lvHZH+V+CuLeRZG8V/RoByjx4Bf7tN79ZZkOUfqqTvs3MHboSYByNkEXSyZainRFVjG
0chkVQr9rmW3pKi/byOyOeJ0Ii4nWKfGDGHS8WBF0gFphUltYDm+Lyg/z9VUDXeuG0r3Ga1812cm
58+vxFHeNwM7gxF7u5b6SHFr02lVM+ySY3qIr6UZg4PmjPikxDa/O2AJAy7tg7mBap6f9OGDzi0d
qqzr2RUl+r+U5RDm850Fp8rHkmCvzU3KD5HmzuFedKmK+QGWD0Rt7vQNq6sg7XDXLMiid/m+No9H
bc+l4p+XPE3Dz+bEgglld8Se4qr6otbaWCwKes2Z5iqFxJmz2xQsRRF/Y5Shp9QlZitJ521Z0a+C
Bw/taGToVlkP9+hnvgdaygFqlS7aWK9ZEEGkM22QQJXlpXseRtnFJPfyjvPruyMUxQDnAX5rAGW2
I3S8xKXRywr5G/RTB/VjkJrE+2IBwQlrOVTQxmwJ4nD8UfSs019fdpyb4qi3LUBwQKKOn/pFIqUo
LRVRU2b/1Ww9j4sFhAP+FkgE7RYgcEXZ9wvc45qK+ctuYJFe3d5W/YWpdmaYlwlgXh2FMSdBbgjP
cVdfctIEgUBhQxDmcusTb9J22KfRBbzgbrBRGwaAw8CfP59sfX5JSGVs7vt6X0ma+fT8XilRm0xx
gUlkhFmd/ixC8rTqAg/K10cw2HfqLUd7Zmp6baBXnU0MwuR+EtY4t33cxy1c4eZT1JL8HtDTM/qj
HTJ5wDMz7b2KhAOGA91sN2afbGqC5NQELw2fYhwP29QQdFCDGWVN5C4z5qY5rCkLzOGHW5Q94S0H
WI/rQe2v0OI8Tlvv2aEAbCxeSd99Z66sJj+CbdAwvU37Fu5j2YZjs6qjxTyRrMB9UzoWcjmiJZSD
bE6U4SIBXUPN/YDr2jdHRuFbfar39If2pLeEDFk+Tc4LU4tLzNQ/SFVGPIg2Sko7HUyWdrEf+hMr
1fQM0+JvRmHeQM/LNDQ+EyVDK2kFsaXHRZvTSbilIZUMJjogdO347Pp7kXqHCif3DEHs2NxWxwGJ
XAhSMfWmmpBLuCSreNAAOkp865fb9y01URnskWESIMOeuinz5PM9KdOmB8gljMnQiJr17inv8fAE
/3kn7Re5rRlAcHU377n8VS6dlPuaflLHD14TWXg0t7VnYp3G5DAqZ3KcS4QTK4Mmi9jXyjOl2S49
zzTZgJ54Q0mWr5U6OAYa0wUkVz0TY5EiKIaMxYxh1UedlKo28QZgH2mlIPOxNVcqTVsVJ4lrrvnN
DP9U+t9/kIBXEdPD44awExjrTiO5cC9VquwhmSXqCd1C0TsHUWZDWiDAATryVGUo20npgHM87Cha
Kv/hOqDdDc5Cc64suy63Yp1DPcvn/ydEXl/ug41cMAO+s8Xs5C6/2pACiYydqfAefllc7pvp9Gb5
3UB0ShlFxlYX4e16AGShAAxpT+HH/CGE046+dPbBbJ95T62slHHehqgL8nBONE+OrzgLzU5Alu8n
N9iIDQ9nYU5mkAQju/Yy/UtV8FpEfM8x55BvPBLeDw2mWLItEOzUAatuPtMY/98rK0Ky6hIeS9cC
TAK4FdA3Y45lnS5FVZ/ABVosLp49vsSMnq0eh5jZ67MeNcJqoh5+r75Gnwd51FxXuUPmbEreov8S
WsUEuRHGc0oWIqVGaSxF4bcTtfYmBx682LtzO1kHJ9n8xrmM+6WQrekiuI4XC9sAX8JPy89NV8Et
HNJInbAZLvXAiZCKvAxModXgYh9/8m2wT0PeOLSo9YrQ86YOYD2DVMX20cLissdMPdTSYtt4RLRl
yI6AnenHrAWcQTLTitJkAH9uArNgODDYBTHCag7DA0Qv3ZrhuPDzsuyDX7DgeYiNA/k1PIsIFAtG
6YN/dPl61UWgceRMP6QkeIhQrPuDVP/o3yNx0hYQo52y3EkhgS0sMEKHMevjp6Q0dzWKetyZqhnY
oR7+NMfBxyGjG9D+di5SSBgK7kUVBy/oT54cCVfxmS0DMSmzP7DnIxNknPscEdiS88IsIqnZg9l9
D+uVQEWrUsjFZuMwrDlUl69adcGsXGjxu+DR81bUtD1IcAJJdLqVkJdIM6qbshYqqsQOKgTCZkPM
KLPjC4ejARveWinxWAya2wTt9pU/9K0nvAv+Ta7KPszHi2WYz/aynblGncvnLXdmeM4mpb/fUxJk
kmYzlfxyPVFo5N1duVVc1EwwxK0qhmOwty1RG0yu3nNVHxcXULjisC/jGfh9ysMToM/QdMthVhiE
1qX0mEPJtx865vxrdE8AelykHLMhWtyxvcyZjhtWkERUbTpRxoDQdp+yVVD+EwipTMStLA0KsS6V
30ZUOEOUUYZ36GQ3nHmoKJCppMAki+vn6L5fbKuTzh32yEQFvCoU4YYa4hkNexxaSgseL99dmRwd
PRmuITdrgYWK9pW9f8ZbB7V6tzH+3U430cGmG+H4Lbjtl/uJ6b+r54YfOm7EJoumJDdjbMkpqN9R
6pjn0mDkV75Q4mdT7aToyfsf6jSlcljJec66xHWQTUNlQP9jgZ4cL8Bsf6/KIK5KvNIKDC8lVOM+
2ECu2o4nonc1Nwr1XN+HQzBLnvXK3B/drJKVKv4GpMjJUVkzu6hOintVbtZxEp6G0U/3qKX0ZyK+
c24JRooWRSG51m/h/oSli3p8dPB/LKjoLhD97lQdtxHEuoFoVRh95beVEO5rh9DQmf9jmvUrSByD
jla9EcV6Z32L2JK/BoWkDfx5XrasgvNVErOnn6OQZ358spOjQzfuvQiaQgsASY4Ysy8wjNDakigS
oCZPV7lXgLieS5tPzsocV8Pbjm8qPL6K+A6DnxEtCXRN7hKvK7zjhzNW6mITs370PvynoBPjliqt
n03OhTk5rGNVgaIehsrxtYloDAJzZtkpQi3iVsduKELCki0o45DShxmCA5VXa/qqnk7WVS2tL0WK
V24aunoHs/mD8VZBsi1E6N2Okh19J4Zp8Nsl8TgF0qgqnMJs9pFy+3BGoX/HLudfak+NeWq29vh1
QRqk1Qop2wDkCNcBvy+WdF5Ml1Z+JEacbUDNvG7YfXHhp88EOpglzZtPRCYkNHLtrz7PX8ECSd21
6I8+yRwPvc0FnutwT0CWR17SSsWHpFRp9ptw1G/3/mmlcUFrnGduXWDzb36BdcM0zdtPzwqxwTJ7
GNYr/mOd/drFDmTSt7ahYFTTXHHLAirB1bnNHdK1cGzMjjySU0AxfVSQeXIGZsGayvq5k/Db8YOm
UO2ASHlCyoeK9haFWSBlBAEGl8GegsiKTpVMCQ7vwYk88fzms6e44WnmUrlf9hMn8yd/a9kt7h+p
VwHbGrMit7tqd+A77eg4Oj/HeEAPuZdIqGNdm+UHhHoet1y8RrqvsfWoNw78MrrZYzY0boN6o9k5
9AcSm6XVYUg4BtTfrEY4eEp7A1z3FcKrFwjzc1jrKUW4Z+verxz6nO94cBPo+4/voS2VnFeB5n72
JeGQyc6ITYofQJUtEZ9ICHMRVWt9Fy0o3NmQLnEDgRGO9BNFMamC4f1oRo4l9IzEbAf/FpjBGUP5
3LSF+lyKxC8r9DPtpTddMJznx1qQ3lN+UYWshsxyrogkjwGhFtmKWVtbPMPSrSL9m1FsOg2OS7Bm
FQXpPq1jQdC0qFds0zJhlS6jdiZWBkn67ow7sOmh5aajbZtpiOlL7w8Ks59DKhmvIWv54rZWCW8Y
gfxpk+irHdMPXaKbHMt9vXtg7crhyMTvPc5ppOYT7YpxSx7UBn+JNwbX5JsbNoghaheSyp26CqBO
SbFx5dX5Lvot28y08HsSKPDztqBktSg1Y2hCSRy18rMtYq/JzLCyyNiv8QdWjDX5mLrw7bLXr6XH
J+WC2EmiwPzGQms4ztQjsaK+Qo/bUDAx8Hk2t7VqvlpokG2MaJxqX+/vEcfMfd86Q203iDiqXCb3
jId+qt9Jz/p7iY68v3nDjqBTU9ExF6fhvjWv7dXm04xALCf8Fqio7DN2hSUodyB+2alYid3/Go6y
BI03siAz0yYuyPf8W5HzItNm5Hw9MnA8M0E/z9zSTo9QJLe6YA05Z+ZYIl4x2BzCTMntwR0wIFGd
F5cPiCzqnhHZ4Xip3ns+5pKCy+64188S7LzJQPA6ELBOmIC0jQFHmbeHAXoF3dwwvoQEMDuZWseW
ANAZnC+wSWyCwpa1XXA5m5Nj/BI8t5T9kjwZ4JSbyzjwQHBhOjH7MHa3qSd2Ijr8Yc4oCpPc6dz2
/ESNRw4KVmrr2VDdUi95jtWPmz3BXMu91O8qcc67I207V2W4HXMhQS4LI7Kk8/y3DjCu0enBENVf
u0G0BDIYdB8wZX4qLDBBGbWJtgn9bF6K/W71F9AYKEXG1WNZhgs7O99QLWuijzAzZyldj93OcQf6
EmRdsnyoEG1SVaWLDLAqoNaAKs4JjYPA+v8zqAmbv7gjD0hJrJ0kwNbaj4lHDDh7syzU3Y29MANf
MDHhISLql7H8h8Pe7rfcfslZQIvvwOLL20iR6ojmaAfKfp+2P74AW885LaiwK5LfUlGQjHpiO0Al
dsWN6ibacNYIe8+HpNE94M3V8BMAMQeLy3c4BZ42FhlsteaUit6CdkfKNeNXIn3w9ULAYTlElmep
DvPa/4yyi2lJYJwKZMimFDlLRX5Dj8zoYE+U96LuTVAv5jAbuio3y7CQ30GAPpofH6xzzNFORy5m
20Z8f0FF/wb+NhtiEqk3pee1tUaNjzcmpEnywd67B01YaX4V0rt5G11OtGqemVyz2JmvAes92Uy9
CKrYz/NNs7ei/e3snVRN+EtKzBuLVkj5HPHUZjFLlDmjLfDVAJlcajMa6Qa2o/7UtaeETTscWxzD
pz7E42ps0crvdIQ5FhQcQppFCT/4OP1Ce7BK2gNvcIj9w36i+LtB6eF0hfpnAaUD1ugRsCjDHIlf
YJ0QK7qnCgPNqg3IONO1JG+IzXL/OmQdqJEM4ufnL0uYoOhSHPiEMAEJDAr5hwWhQeze3sFS2q2/
Q80Pqp6L8spqPV7mOgpynYCjXu/KRSARG8QmkVcWD0Qc8xaguskNxQnpQDsVeBhe3amSLqxEs29l
pL1YIwG2ZYxHicuh4hSoEhYQmngn+Bf7Cb7UbVbn6AUpghvI2/EWS041Tj+k80U2htQyVfb8af/T
jGPHOl1LBcU3zvvuomniTNwpoP8RlOQaq3YG+2TYgD6bnyp40kfUp9Uf5R1L834mJDiIs+bWJRBn
kETjtRn25Oo2WR6Vf3SZjQe4+goHLexerz8hIPKGJ4uxnoLBXHRQSE5j1zjUVekBXEBPVidEh3cp
poseuDF9kOU4tKt2rD9wa+OLPeTS3eQgdVAfr9/wlRMzzKmLc+5n+8dD6AW3HFtEKLginI9T3WN/
eLuBK6vZt7U77KBMgnSEOccd5N7NiBR6BY27Nm5fVD2+g13WWgsnQdOTk7ax8qqfIWMmezE4u6VJ
paYa5Dzt3Mj6oCjv2Anyv6ioIdXWBXCuiYpPAFxwAeMxQ/3pEkW332t93PFQrD1lMU2/Y7mptcZt
HpJTmTzn811dfCXW377CZBVwYi3vYieJhUUF/ZmgapfTxWgpd0TekmhJQbu5JhMg5PNzChMp8Gcr
IWJBMt3Xa/nXgpOWtFw/YaAhuUnElDc5UydEfA2xiLmZpwoeNtbxpptSsKuIpJSjwkyXnE0YOfgV
npSq6o+n6NVYnv3B0RfxbkOJ+hqECRDOBqmQoG+W3dyF4+0uEglWethlHrQe6sgycDZc+od6g6U/
/LGv/RwKL4UNBHJpVcfx2GPqxb3uSjAx4PT6YCgdJyWjy+AHTgheznXQTKXUl5+0bWMAzgziL5rb
SlzlQuiL4JWgBAPsFHy64LlzWaTRlANYCMeNIYRYRTkuMpH88VooC51vaxYlCDCUZtgsWoat5TW1
F9tI3gSgQZauJxkNHWTpyKK4Q/Ky8cvq2pVHkWdbtlW7SGT9wzccByUpqa262OBfEzPJ4FYjyzqp
o4uKTANl1uJhn/pmFT46AzpmPjTKC85zouNEIju0XSceFVKOrES6K2o1Qi8Ay4rZ0x4p21vXuJw+
9TqgS7UNxcGOcVhqvx/TRhlSwUfyahkJPjx+dHAZcqElEE1hrtxgV3Pt9n/WlQSc/fTJkCXWF6h+
Rr4wPHIUyB5zMl/VayPTiowY9sH1sPaaHn28sw81ALEQRXnbfTPmFJrzVWKDeI8axWiDvn/WSzI7
Vs5rHDTCLK8VaTYfCB2goxAkxnBcJEnka9naRRBd+adfcdjG8EhRC0P77Xr65Wz8PotT3qF2V806
rgPDjR+y/1f9Q6w0CU/4uw6E/ku87a4XoexI356YpNifVTF2lYQfFRfbEvIOFY2fYoCc8f6Hk0Ym
ZN/AK+jUr4tIcbaDhkg7+CGOoogwImbfU6ofD9SuqzMMnp57VNDmQry33QhodFmrmHoKXDXe/nsT
qwINY+BwTat3uo32+UNxhdJDknjJxiGMdP6Pt+pbqU+ym33CQS0WNB2EONN2q/IgezNgRI0tXzN6
54ed3/AnKJ42I+EIFy9dOkdnFoDdUDdbJnHSwzUrG8LupFq1C6Mp+v+p8S5q0bsdC8KGI+T8rFkz
RBnCFxE+Gp0MnpkwK4/g++7bL0ijMg4q/O/81Gh+2MO2iMb/6IUWPy48RKv3ck1wYX3g6zai/z+p
Ocpb7SD0OYRbEGdZepXhS5DU53H6xq7B1KHOwJ0DFx36DTMfSMdgNYp74ggJeN6t2sGowx3o6no7
EgUbi98uJkwbn3FXcrEV8Snj7X4qXGBj56D/n4f4AlFZCpSnaw6SeSK7qAZhpkZEfl3uPnqFSv/a
TKZLKRtV+bHFCxssJWfEwVk6nreqK+cEqO+sZDkXl6h7N0aWDi7RHHsbchJiK/ts+NQ/oeXJK5O/
K//PUGzOTJFCGlW0pXC0nGOVPtMWrUqG4Oxc6sl3m5JncK8yKR0T6LGo533HJxMvV6QWGgX8eyde
s1b+Ug12WjiqCmuPSm2CLYIIV8/84wo68V8CtZyfGdyeodNJhdZClAv/2k4F2WKx2+mU2saqX9CB
wWD1H6zf2KufVmmY7qSjqQ9l6JYdyDRvB9uC1xQhRL+Bmt1LXHOxxxyK9z6Q6vqHWdHOTxOP+PxI
VnoOgZDdPB90jyBlq1HlCuyJb63bRbGr0sndzp3XOq/K4W5F7qxggB0E08+yoBGNaNEtd3O0v0SG
AsCIUqL+fvkUBaBCBRneT6o9CV6MKaGHsI6EyalHju4ifrYtyQopjmoX1dwocCrVw96zGyj02MKW
Gq3FbR85hSYThFk8CxohXGnDniYVsXOracpHAX3Dtfzm9U35BWWUmbrT6Ynlx/KI79WjWnbkJZh3
SzpOZSEdxY8xILg5GnHUoCU+gKHe3ucp3Kuo7ZugXgbLqrPAoCEFl9CUJn+GUerknepHtww64d1o
PFR+kUutzIikU36RLc5Ro6CsmDZEsq2F30rao6I4ei02P21lu9pK9w+/RHykRrkj6C99RnDwAtD2
xX+ElKQcUfqFDxuQjpH1Vyzoew6suNVCpmwDHUVNjfavH0SsJ8T0nQL3e8+sIFPfqC7nQU8QedR2
91/wYX5CnvQUifEsnQ+fFp5DNEPiOynyyuzq0g0DOceo3+JUWm17mpr14EpWYJiqvDzMVrM3oqr4
yAHQP6R5zYPqxj0ARr2JPnPuXfpA9YlzpC5TjznP+qZk4Ei0z+g1tofVY4nEnpDH7FneVPVJqb5u
Nicf7i44/zkcsIOMI88nnyL5rCdGZFO2RV7EGBaL8KCFBURC2D0HEvNXP0WWrF027ZmrAlT7a7nu
Lngkq6pHYgceHl5A2hT031H8YSXpkHEVjclrerAzAu+0M+e2RrT0GnlZxwudImYiW4kYRHNaKWS5
+xbmAWUxI7xRsaW1NsLDCabrewgRQrm8zdCP7bBp83IiyuFN/VUot9LEzr0Ij4Czlu9K4fpw+67B
hPvrMNkcKxv73z8oUczXzOshh1iwxYsuwhnxhQ5zk+tJCkydbEvBaxDAVYcTt4dMMkjdBYHsZ9VP
D/GfwuWrJRKRGFtHp9MSFGagEYHMPZUXSSQsH3Rt1/8cU1Sr6Ksx7q0GYdQKbIHj0FY/SDXdoP7a
l6P0XgYjBAHPJoV7BLrbGwaJrexCz1nSzH7PfMolMBR94+bkFwCqVUYDCDJfUWRjwvsuToP6Pc+6
pUzJL0nI69nEyjlOxNoGuXu+covVwAR84eEQ654kwktfVFNXhRdZaN1HKxVoD6IDkm6gQ6bkgh3c
Du+ND1m6EMIi7d7SoD+0z3GaZMJ46GaN9kDj884RJHgJ7cu/qsiPy/cTvBtTg5yJcfsQiauRInmg
AA16LKGCGaxt3Bm4VklOH6CxYjvgDiUNmcaAUgBjWgb+cNGeMoMJ9b8TVamIDvy4jHzC3T0GnCJ1
EAYsoOKgGuvbKPYEw80oFF9jnbQOKZxsM2syKysH8SbLQsrgvzUAG+EsTmhz7wmuFyMNn6m1aSjd
5taTEBM9pTswTcpEdZG98IemJ2H7qAnhhzD0eSK0IMjWsrjhZAhfjywx+2busrivCDBsvSNrSLot
4T6ssH/RtTpg246ughGc0XPyU166to7G4KI6gcuUee8r6NTz9JX0MN3+vbkxUT8pRCjp7+Fzu7vS
DiDLfV7x6Vi4JZgXOSQIsxGOt1ycsqMyTx8zYYeIVr0Vfh3WdvDSIVtwL+91FWkH0ODeXAfX6s2w
tciBpBIhLGiaXSa8xyS2Bhowq+g/Ej/AU0Kw8fCPz+BRdGfD+EVTaUW9ZvTH/nHaKPpPqgr3XL5V
JftRLptMlvaUgeCpscIQ+UuV5pCbAc9Ot3EoWlgkrg5ozRCaq9lNvu+1tKXRMOkC8tvkE7PTocAI
WlYDa+9D2pObYoTNZtqMQ0rfbApp2ZCchcxBZLrSlrkhyj14qMbUWIn3vWTAAlnARV/HeLYpLqTd
UmzW2zjuSgg6uaMW83pOKyfngIivzn0x4Z4ZgWR5UmaP761XcXgjMSdv5ARD4G4REsbzG5kJEhOI
a6nbjom48T2DO53OAnVDeAqAdzZICwpFFEyMmZpeARLBwF84khE4TV+FQ79PgjObDNJeVQTj+/7C
1GGV3l9xl5tAu+fr6j3CgudlGFz9bH2ezC84bTa8IBPwPwVgkE+p1b0K768mz77asN+fBELuCeRu
oMwn5wvDORXqcMkIghx82MZYLXKBd+lwksnEYbOX1yuKof9rPMvlJpbsx+pJq2gFOzyn3k0Hh6Tv
IgC7WMJyB9ZyE4j0WjLr4i3spzDTfh4+lNOrcIgI1b0aF3mIBz8IPibCd10xKo15etnJiIMWgVgf
sDWuZtajMBtnTg/9gkkBEQuOhCZGV3i4xjoaBH9UzOwDoBynF1QdFrfNU3lFEcCjWUAyeAa7EQIj
g8T6YkufgZR5s5Ch4EzPm9Wc7tb2/MdTsGeCSovcUUQsAo4ZKUvvMYt6x20Km36lE2hsdRIORHUR
zB56WEvKo+NdMf0BxGkugc3sgKYBJo6XOjDPCgA9ZSoaR53Iz77rpDMVJFxEi2Gn/fYPDLcnfWfC
y3KnneK645zvY/cEm9XPVNPOXQRyOP951/2Im1/Ld9o+A2YgqxUZb2vnrZKgM3xZmh/RxaW4EmXP
F+kJwXgClCCBTYtjrfrc+loPHNyniqb8ncSb1Bq2Xc54+fJuKP+pJeKNkKya1sm8+EPdM/HgwGws
IrZ7c5xm+C2C061pvABsfxKTvxdr7vTaRwNCebNDXjBnOVjfvWdidGssIjPR3sQmtbcYsHhyQ2NA
t+iy6b+BY2zXxeKjfF9bekNdQ/T0VjqNHJf+uyKuvnhdr+mpCe96hHLVDSNSqKbLJXI82Kda6Dx9
41U0kf1F3nepFGZznnSXRJ5y/ks8jMNmvfJ8667ZwGYZ4lVnaj2+lxPtRLJYJBP14rdFvNBRX22P
7Iqs1oQ6ZlD+Dor9+HECsBtza59Wj80MzNMtsHbNCRb1jfiv/isyxZ0DaZTrrEvE2LeMe8NjkxrO
TbOOSF6fuOZwJOGm0ZOruj9cuRrPOJU+347xGfNPzICn5A2lZfdImo9MCAY5EIlt2fE+flLk2BAy
V9IpPrmoqsxjw2/+iSt6m35iOKApxq4YGSF9/du8u0wh2vWaQYu+09OF24HU8B8EHdhEaBMaXX1s
CaR5VEzVweveLPjFZFTr9jHCudLCpkZZHzllF9PyZuMBiVUoj+wO/TQXZEyre7SGmKyRGQvXGeBA
dsij5qJsFwAZWAUCG29vjWbsJCvxh5Jog0K7OlRInPDzSf5+WZZQ33XZ+OHt3sQs6bIpttfebi4L
Coyf8/7pcc4rbaxrl/mSUOoO+NySWa9KfdN8rY0uXCYRwIpJ23TeKOd9eeDTz5k5F1kUF4FsQRyv
ELCoyRENiW/fdfmWC0O+eliBNMtcCVO8WTaK9IluTn66H0Ql6BYB1itECfe+SMM+wiLfFO7UXCmw
UuOHozN4yhC7yhBFYjaWoP+S0vbfy5D7RC+u3z5t8TDWCI58x8wO3pTdMcdjvKWqIOwl2aBpnTSf
wNVruGEKd6nM6YQHmeJAwKrU/uXbDOlMsufrnLIzz43Coi6qg04P9tPZGUTOwh2U+phHP1/XiJaD
d9qK5WcNVAvSjZ+MqSeSTAeEjp9DW29HebfH4taOrnVez4gT4E15mGF+/E9kMuQ28msrXtE7mlYl
iOSjULS9UWworR+n7ZQ9Ux5Ex8E8RlakB+cIIU/xrpyG9Vct1QJdyxvrwiL3bM1AnnwBZuyTQesb
HyD8nLwCOoxwF/b4NzLVVAyCo/BrZwtetLgxb5Xj9yMKEKoMzv4jrD2Z+PvdxsLRlItFb/MmXIJv
DSsePZ7EvjvtR2mCUT6ldehIGJvpApSvpt6xWJSRY58PKjHiuNQivYyb3bYqbdPkGoWrDo7pwf1z
8iMArlcL3jMVspVYIPGSh9pTTm6mexBCxtzY7EvZn2M7b9w2I9wxUYklqNE+m/KM4Xbe4JVQe+XY
FGq+eBVHcT8cWlPQEFR88Zg57B1YKnmKPQLmA36/ciOG4nI0TwzpgYk0LqxTKJSReXN3y48h630w
GR/SXYL+4LeeqwU0P3qgrgo/8rzHjVIXIABnpN/YMM2XOp16GzLuI8XIJQm5a7Bpy8GY+jABFbH7
wl5jPCrwdq6xqTxbwrQpf2gu2MF2Qht25IV9Mmdu57wcQZ7nELjZTGVkccT5mngEiimJTCgRhZ2K
0auOvS0zkVa5SUphpSGs/mgYTla76flcZrkrLcqn6V1Wy1Pm2CstTBmn+9rF+5wFpu47xvCNeJVN
GvHRbxchIh/ghsbNajIYsQaCmQ7u55u2VuJA/24Vwg5ofKBcIqqIQol6fbOgt191uSHTHZ+gnUil
xH4ugGscpsR6SR72BU8ghPNUNyUNDWTmQZ81rM0wauB7ymQP++qPaN9lxNBtYYi73/oSWx4pd9HM
jnSVQSM8i41lznT8JMOIo6vqFRzNgV72wrtxSDib3Y6cfpw+qhnWiG16xAVQXkFTyOuq+u7BtnYO
lbDeyGwfHQPfoWtR6YWQrQbnEtzzOSHIYY11J4kgFqZxfaWfwF584bZfNE/ri+mQa/7INBqQFymz
x7wGuB3sv5rDWjwR4gyN8ZAhywur3dmiBKwSNnfQd8jK0kEVrY2+yAVIiYQCpYRd0XXN0Lx3IRTX
RLGIvIi3nnPM/98P2OZznux+gSjxzk+48BZKlZKfrkUpmZCEOdGaZ37cwZTEGWYX1vhuOsdVcOtT
i6zQAuJ7JAfRAEziVVGFZ0NPMtP/0Svu22YHygbwk2JtZhHDzzcksEZKpnFmHTauswySVqXpgmPS
5Ztn6+4gJZMtem2H+kARqtsyiHmuwTmNLB0pMfc9y39EBdETHW6WbSCHe4QFoO8kx6TZ4gIC1TDo
UKamrO/mJXZW1wtEL1OsnWfcNYZA6wIiZT5l0iVXZ/arTuWsfpG8CxYqLHQblG0WL6pktALE9C7o
95dFG7qeAQVraCBLA1ZRgu+C7HCzOK0kCQb51d+14srzdlQ1wve6fUFHfLZd9rL8SoeReq2I3bz6
qlMo7RmpTWBiY+ObgLDOgZ7m1iksvdnsxA64bGaHhPWxVoK0K3se+NmeXBowJYXMXCZQ2iEKxeXS
SelfYGeVAsrUjs1gN+f5+5kYwNdTKL6SO9zJQyr0GIClOpMP2fzXsU9g7uqZX9WjnnPUZq7YpPkG
EKKNyjoKeO1tYAchvVVP0jUPtVaPjZvOxYqUDkIOrgyV93Rn/yKdf1JEvIodEKbwnCQkLtO9dasw
9Gy659pxi1NajdoNJMYMu1M2TYnC8xEGaaVP6+OrBU3HKhdy5atnCYjBT6flYu9q9iV10qM2LjWe
/mL9jEHH+aCaO400YZVk/Q2m0w/+1txmPB+XTS7dslgtOAB0Ko5Q3rdMjSeppHjsNA4CsQ/FFlHi
8m1bVRrGm8mqBZomukDhRUK8BU8hU0+74qao+HcuueK46otidBxAM3Y+URMsTGIF+ZsxpKvz93yG
onucPjfpbKtvzejEQoJRG6ryV0KHvf1SYUXAdxho8ruXmuIm9QnvZk0tiNtNrTxMa1XYKYO3svin
915Kj50LsSghSEjGTDWyG218M85X9a2S6xW/SMfrt86nwYKiyn0gWVRFXPJQgXYWTHrs0XzLPN/S
cI50DuNfMCYj5lFGPL23Eo57nn++93YKH2rAWNugR7ude/ss/DjEPVQBA9wX7uTagGGfG60mq5Ti
jQzZd6ljsk4DeI01ZjsYIN4ElvPZhklcJPzJSVdGGVsXPiQWNPtHaMbmksbZ01LYYxpSUjurmjbo
Upz1VanUxcYpenhTm6rskIlOt8OaSJ9tGoGqPxLxVwYPIcpA1leQIFlEdOIpV7dS2QvS9SkpRoHb
G2P7g3FIsxQFyFvfhD6cpo1APlf3X+NamaRdXwJvvvquzhAL/biaHJxEAWZi2mItJw+SWATgTchF
b+RBBJ3fC63pumuXuSRXabA7nDMPSCYxf05Ahr7foKb2zlp0OfrNWBIuAlh60i77WpPspxupGUfM
7VhZXLQISIMag0mTr4DcnM7Zn3ump0t/LpV6jzV4qlEoUDNo8kbvTolY51LYRI6f+w29dxdrBtxA
ttNmdTGvF2+hipfWgdf3dZ1lq6iA52GLilwnkb/HUoQA6qhdCz0P74OPYLk/5lOVPyfXMuSzj6fU
3UCuSAZO9uSisydLKD7V45XmQ1v5Mhrm6pLN/GRtqQRH5iXZek9pNyYWd3BPCa/U/+9ohjMKM1NF
x+4X7Km0xvmgTM33aTLeWVC4pUNo+nmkY0RIDPzewer3gfNQ+yBCeXHzfBvXdJVwqy6MWoFZODou
3BUodLtUamHDIOwuD0i8/UjOEScIfQAjc6AeT/ncSCh2f4ugJOU6EElxyVh2BhFU+Afh/YSiXdaW
21a6WkvU5NSTA1ZhkZlu0hk5QtAW8+hW4GV/muOzrxjksNcLONYGxuRBStzFIESbJvHZ16QmASNx
Vb9yqdBsD0J+D7mfiJsWxytRdVcLQ8dAcOKSbVj0UZRn/iR5B6qZt6TKfm8XKC3Qdfh9pTbdtuPw
BxX8jWaRQMUDRK65wjKJ5FrzMqbHSXhOBI0PWl6M06oe1d7ciVsdNFiQBF6GOX7hTaA/EtqNXL/p
lbWNBAFjw/z9dTKJ+rE2ChA3uZIROGY4KASCV2hJ3+Sojktuqu3U5mjITt0Z7GL6z/iQZQGBBfB5
snpq7NXXaAYHm2hRDRX41GzJH/nvHRQSY2fvgWokyF9uf0lkHYI4SqGowcX2s9dsL0oJutfwAFmT
39qmcx7TW5nPaRqnvJ8tRqBDSqFnvHDI2yPJtER+8to76oUHq37UgEVg1uMS1S5O1wLLTs1Vf82B
V5NcU/O8PRbgS5rptfFEf9CxIgsBxtiZB0wTv91RejejLwO4g2Hy/YgFmQgV3+pMMScll5Ca/kW2
FVAwMOZ+peigU87bjqpfnudPKIBC07Tknmoow0vaWbKVWHa5gJviRFh6BQTPDn0wOlytH26WlAgG
Q3AsxfxMy79Df582Oi+OgsInm29pcOb3tN1tF4Al4oB2ORhqdEWj3JQ0PLwsgzNUx19FhFsWTPku
mP/GMFuFJr/OAZTLf0hg5EQDLEi7IVVYMHEE4HdgyDUlqiCEDDX8N051eziLubafY+dyue+MqF9/
n45F1QgbwYAiH914Kr8DPC+qwPo3Zzr2uTx6KOlSrxfEi3pKgCckvrrFRMpLS9RmlYMH69+HUUDU
9s4v1T8dFHVvEOvdhXt+krVSdsmTMWRessQ6hCWxrnBg4seVu7dXMgUNKpQBrpOa7ribLR7ANuoG
/w79o/2Qhh1gtJ/7BjLXcQMyGYJYNvpOc9IKhwFtYgwVHkwjZYzsqBXr4WiaycOJCKRHuUZDaVF3
dF1VkJ77S3r2mfpB1OKKOciszhp0F9u4ITsIXXfzfhuFRrZmaoD0wDEYtYtTHO8F2uYIsiRzMhKI
ktwFUS7qkOuRUwnh89nuB5TKBJJSpuYebhbGVmSFx05pYiyozNx2t3KjrpXYkArcM9otaRauJxav
eu6FQ3WhuD71VYzCdOcnqyUeABgdpTt9KU6Blc0vR1xozkEwi97BdDTeZ9GIgYeNjKfUKOsvRTgO
z5I7Iw5QR/72Tj9BiKAtFaDbSYW8mmIlU3Xulfzo5RbIhYJPIvvCFRBFqgT0OaFlcug4wW2irifC
Mb0LTKmZ90WyYBh26EhEYwEQkrBBphKk61xTO14SiAb6P3JGDWpESixIXA7jEq5ctVrlS/O1RJcv
Rs2hfhxA+C+TJMDO9jYfe7FE41S4Uontqn3lXCJWpjnoHNd85d1I9G/kVGSRTdCKlLO/6TCO9QjC
HESXmB5ZQ0YviFVOS9sHK5P7C/E5rRStu+KD/TRybuddhgbANbguBK1q5Gnsq3HvdeK6B4tqnVyC
rFHLD9mSEa/2Jl4wukVfRcFMUdgDXuKQdhnm+QSrED/NGj/BeITRqw5qa77O8nOOTfSW2O7ZzCmS
Jn3LE8LLFGs+psAwope8tIwn4wApFkncjak6N4govyvsu8X8WK+yVkh88vmCwrbdH059zQb5SRi1
tN+Vxf9ot21mBH+y5x705Tex0AAqWkLdeKbM6aSOCWdhaWZ1TJ7d8mbz+Vjh6qfS0wOI7oJNJLkg
TcIpDrXiUrRY8Z5L7qfb5ji5+14BxK/HsC2/B9e22/g5cd2ZGmf4H0jrAqC7fl7sWcVS6feL59ct
wtt+itXhFCogwqd1HNtFhmYQOpnCoqSXpIOe1XW5ckeKnMBMX8f4TTlEaVzVjC1iBah7aocraQD8
0teasRjY0eCTbqT2wQP4uUCWm7azM8xPyGsHG6+zicbFPpVCNTLa5mEwip5Dhf7ZEH4MtB/5LK/R
Lil9Yxp6Bj1CKc+NflGnwBe1JFWGb2UUAr1y+/nriLHkuKHKL8siABtfXLYGtY9Of65WRdusZUV7
nAe/Hp2tUnpbi8r6IB3+X1vgyu2kK8Hm7JTeAT40w51eQJNM8vxIsRBVZmBEnfAEuMb0FHDVD1Gz
q3cZUklOCA/C0/xGeTgA4Wd3GvbaMvRGInVrifmc5KVJIOJw+Oaoa/6dg2NJwgvVL42RkFi6RGwf
OK93HcDz5nQBiT0X6TPYeyMWy+XtTZy0TeytVYVqVLdRboTuHlDHgFlmPWRZr5Z6mcIFUOk6/dL5
4six/3koXjd2mTfigPdMqhj2/aIBTfeVtHrMHK9Gg5d3tN2wAQyOIzADL63zM+B6FwlntdBILYpG
V1tAP1LUZ1syCu7lPL/E89V/3Y1pZ0bBjS8utrVicdDQEc/aKqkfmR7+KkQUbDsTXUUFt7lVY1ml
taeZkPaa39KHlrgC5DvQrArvfiPOF37+3xK/VUP0IkLO6IWIu+qPuqcWdbboL6x3TEVfGbBmjjXA
8TAApJwyJwMkXmCirOkwmbyguAopd/QjOhmQ2oeUOROcGY1LsNSjbiAUONslXzjWlifIqIh+RR+c
fDYO/IBg4906pVeNi1J3Us+7s9NA6AXIAR1WXSYzsJc6FUga5kExVrljAhKqpDbuD2qbNY609mXF
taXqfxwnihpV/a1AkvuGDeA3YhqC83LdJOlquPcAhM3P7rMzYtJMKx9vuQozoxwPpoP6HFrv1Aqa
Xdmn76GjTbfTCifQN/YUceJIKVJT9kYNF/ClhRcs9DloOofzrFMsk8liHDG7u5+6NNED2hTMfbs0
/9qzdKwulVQP3FkiGyGA+sPx6z5omSLJGz2NRe9iKxiysQPe6SNfANKpXHiQqaQ+dgxdZP9dfCSs
jbGKUyYl9iU4A+FIAbI7eJci/Mo92eIb2ZQEQE/iGQIamobhaydMWwOI6ZgnnpFWBLvPMJ2PjUon
cIaAUllvaPY27Jxe3WJgGMN5pPkyvxbPqIKHFMESayt4k2rCY5MDAsslKV6AF2l6RYLvk5iakr/H
tD+jMxa3k8m9NhfUlpulT6DSEFtSnfe+OhkRv2jy10RerZIHinX7VR1rTkHl1eYYy4pfb9hQwP3Y
W8DKFjqJHj4hj5MeLpgV9j6mSzFyx5hZY1Rg0dHPd5VnvuOYIvU6AEG2qdjj/w7HrRMQva81KmkT
/U0cUVR2qljRgAjiVNgfOm8QbaDf4NE2w/nPOG+MqlIEOs6fJwOdhXB7XR7WzaHktBHPKNlcOQ2w
iIfRlDOmhCgFOkvEbJCNYpjF+dvfSRYfLfesb7z2X+wVCUT2fak52UtUzUTd9czWG6nSn+V7dviL
8oDDAMg357LCktm5Exh2RwjLD8m3NdLBykj3tNo4/8kHoA0mLOQwAEjxOEPMQ0nP/OMliYdxiGnT
3Ulj6KIpJvkHuo55sTl3q/FYgKfQbKSS9fgI/0QA1Gs1FIslcP/pb2m+kEls1HfLIl8WYBk6QsoV
cNVlTReNvYRRnkTrquwiVSsUp4t1oGAAF8qoiQCBqiafM94LaylGEejuo+T9LVoheqv1POwJ9lRW
Gf4H0qNuRO8/V+QEyoPMr2WPnkfHm+axftrH9g+4+S0D7+Js1q9VksiblwbrIKN0+n7JndAOExd5
nGkYItrxnpMgydrkI5bBVNiOm5O5ZYuTE4v3dMDmg7NUmETTMv31TMyhK/3zRsYsQUuEvwt7Nk3b
Hg/ni2fcHdJwvDexdopyLXCmkKHlND2UDwa1AEVHssbaW4rlsZQK/t0S0wRjAqom/tQDVCoYwSPh
iCH671BrBAVb7XTfqOqR/UVl+DFnDU+VnJtsUQalqYLif6JH7WpueQ4DgiCO7YFBGxDDBdAnc3GP
+Egxmn50/Xy5O/mVI9KepEClJm8bdOjcgNe8Dow87Gl1Hw9R2KtwsYoqdPlQOZXkVMby9SHremFp
idCg3EAswLbErmDBiE5oHffIP4FD+Hy8yZvwXQ6kQRQn4KyldLP2A3Fs4CaWalNQXAL7FJbOZSdz
ytkdys+kr5ch8iV8vIgmUuY94zaW5UiJwd+1L5D0VAhM/6mC6n10o2qtd5zsGaXNb+uCwn1vr31Q
RBhZecCW7sSnbvEgl/SyQxhL35D0aiMLJlTP5ANFIp4gBXrRAyjeQTXi1fA0Ubr4RcmwQEbvfgCO
TCT6pUZbVtSUTFx5VsLQXvumnWOZsl29o9UFQHw+DgrsrCF5ZUxCQD6Ho5sMXK5FUo8iU0+Qu9cN
2+QhPg76KkLJpYFN+4UrqOlmKQ9lFazhR+hOLOKhuT/3Fk+gsz9SwKhriYcgW4ZCwVRUOwA0AHXF
MKfRTQd8xjX0YKbjBiabnX+KLdW6jOryhUTnXVuJ6O2/pOac1YbzmD/CkrjcfMzhu7TKEtRcy81w
k8JBTHh4hApfAes2CW6LPB1PusuIW/z7mgO1Jtb1HsjzaVUvSHEFSVYmDQMJWMoQj7b0URhanz5S
oKbjB5uyJn/MCyO39oz306a6J5NtxYKcB/0dkct83BoM7QqNU9gwTVLAXPwMh99QpzeMbb+CeTmF
urtX9ITf2+ocETlAq6pdoq6tJB6n1cuQ8d6ChgpFd98F38psMEh57RVfXwbHufJ3YFnUe6/qO9Lk
+UaRUxysRr0WFtQwwTffRsCAWNRLKEl3RqXPGKfh6ltjjQYGxKkV9DrJwy0VsHHa2WaE1TniWwhn
GIv16AwcTvpAOBqUrZhz2UIm4O4Btfl3E8ONeC+ssc3cL8fTruz3a+ZG4K/wtVyHk7MBPzAgqiNT
lweG1KGUT0If/13lK6dYycKByTAwjwMuRs0vRL13ekzV1tvMAiikoBan8HXuvQI1t5EC/wcLFWDm
yJ1e/vEIqbNgoaNdgDXpBpdJAKcm1AnLau/1OJYHj9XdHCuuO7qX2aVq1QAxrksOq/MKSgnsAAB/
ZfMVBs4daYs5NJXtu81ZUQr0MekmsCEHwNzf0sqzOuV1dX3DCJhTPH3o3gih8o40nBvHyy6T25oD
lZ/Sz79z7eu1IWZs/usQmIpDc/P1jdh6if6PjfEbKJohb8e8coYdqA0uBsSUvVzgjWj9m9NVVxAC
iVwxN+yySMBAb/2lRT2Qe3c8rsGSmXgoZgRlHsApyq5ZEsS+7Uss5pel3jj3Vcw8V7rCxe2q5SGS
Ql+veKCIb4sX2thykR6qJuCMTSq8b6zK0UARJeivxXjbdlwr+l3/KcDRGn17mmWhvrriBEMpDoaJ
8JdQ1JHLnsbLQjimHETfHq2ORJYlPhSHN28NtnAEznHcKBZeMJkPj1yBS2VM7kWhJ1zE1PSXNfkw
rwTLIGhTUkHbxRE0cG5l/VO8wz054WbAYPRmNnPC2KxAo9BQ3mfn35Ah/0HzVG/cs14nZIal3g7W
vYV67Z1BTIovVdGBOqdhUIcsMcbriCalsGTZUjEOPVrQwWzmtss4ztB/MOTYR0/edrRx5UsMtDyp
qp4IHVZ314wCO45FbQx7R2NcMCZV3FGKaG3SamMPDtWucxhpmb2NjnmYurgv8V4I4DISoYEXC14q
sWe+vAuBviePq7Y8Sj1rIcflWRbVq2wcKBZ8396jT4CxPLuJnAlL1ofSj/YA4xIwjQsva6f9Uikp
DUzPhY/eFFUiWIAzZiia0co33n7YJfeSxf02qNbE3x9mdVby7DUA0QQL3J1FihuTEexhPZbezhBn
Qb011RYbYuFieAr+h7/W9XdBZQF5hzH0uQBeIMlfP2/76tYj0GDKXkalU/UYgpbpVIz6yb1Upr5x
chzNXZVTZFo6Z6RQ/aByT3jcNF0tvYV9iIzwE0zEO1B0MVqkymnupCHaRDoPVmf09fPftcAgk10v
DKs4G+rRup1xj9F20dm1SNgHxd4+LLArJR1wF7YbYHriXl6CpfoZ29JMvJIecuYkIv9vZfACTkL/
lL+ONgrQ5UgSsO1bocA1E98yWkKuW0iqczdJzUL0JNjnT1G2bvXWH4qqv5/ELja62KnJi0naXPSv
yprkF+glvgqb57FvUnzxh9uFSUQk0Ogj8iH3smUKCIJ4c7ExxCZ3Apuyl4O05cErHW2WGd2q+6gk
Lccbr0Mi6SMDmsbyN58q7gP6rAAsXOYuC1g8ZIV/daD+Lortv5oYgqMNlusFyVhMsvN3Q+F4TndA
KUihBrPM9YYe09GOZRhkZrGZFNrINL7DsIPIOX+GdVJHSW1gIFO5R41ALjXvCBnLX8ueyb8AhtKP
lcXhfp/PGWq1CM6Oz2lHOM6VfEaK7eCR/tFyPKTiQfrrqUSpQW1ifHpFSwAFLCk9wSadgVqeRLsQ
2SNnJW5fxDQHvWO+CRTrY8gOcDPuU1NNwin7SHX2joeYYAopnBIhXeHMIOGv7MnwvtUPkZBB7MVC
YKMaUZ8xGgAb5PH0a2Sj5tzHFpMdC2eu+HxIKHqiHhfP2hd9wBhi0MbWgB74ih0w1LiCPZfjivdK
T0E+XbVaItyqSA/mnA/YDvt+fBRNMsUVY6cOETJekU4Owr3FVUHKMcMBx7bITINvdKH5SW+zcMfF
HUjW76Pq/QSZpLtcsmrd6sV+iu36bCWo+xoMgL1D27pYuax/TnaAMkzvNq2dFd1hEWYs3ApP7nrz
yRLSEXyXzS2tzMRVaYJ1reERfGVwrbJXm7J8zQ1v8OTrNz4L2cUgEvhRwHl9dvIAmgRBiB+azNxo
Y6ouTmq0ff5eNKfT+AyEiDEr6a5zEKsiV0o4GnmMxEXl7i4MrUBKETUyTNYpov757Q28z+63XF7u
lFqnrC2tva58huUbE+QFtt2J1Jdmm1tr8hq4TcMfiK25cemZZzOu7Khta9TyFhJUgwB4owrY7NkV
7wOZy7mqFy5gqYBmUQfK+ADsST7ObZ3Z9jpZLZ7b0LDmHGGjetW1JokP0ioOYpPzlSrvt95dSjWN
l4Uha3rVgfWY2qA4fEFaM17OT/vSj5ew9Ndy6FwEVX2aTHhYFw6LZt0Qi2Dn+nMonu8wa0e12bR+
sFTLnlAc3htrgkiKgXV+guAibblGyeQG3srfQ4CaBquZ9rZwbGjmxRvXpfwoPD7iGExBWyjX0fPk
GKX2Kpn2zaD9exM8et1o+Z4xCMNWv8QsmsV6mwKkfteTvRVJVgyH3J3yOQiD6tUvFrLhBpC8X7f5
548ig8bh2gUminzYA94CWeDJOjcHyriN6NnlgyiqP7yHUGwI3Nov85Tutd6LgzBXMAYXl/ClPzvc
pBvcrX1qyrHEKahb4yQfMySOUUIXnNv4idQRBBGVicEQ/Yt5nDHJ5AdI+iOHs5+EaMQ+cb1WE3cK
Y2PqzPI5pKx8Trnh5I9yTRfPTxHUSHkLqpbphO6aibNI0ZDnWEokKrWzM9GTSCVwurlkd9B/k+BS
/1PFleOVtVE9sUkboIbFNU4c5GwQxNBJqe1RtzF1LYQq0lOdpdnYTnhapC8tLY1ys6yybamMY93O
WMD718mnatxhzX13yo3ms6/tzVF1yrmkikig/t9E2hyPJhCdLy332lYYMl+Vx89R0jzByEwoiN7A
phiA3Xo+MwFtmYZrBZtuQk6KYgaR3Dr0hwCJfUt5fjQB9fOaJZTw+6Mlb7L9zXXy3RQ0s5sK6M0q
o49nrT3VOnMNTGajE1pJw7lEb8IwsviU5OJJbgeSeZNjVGY+u6cAvPDS9m1SEIGAIBmS85Zm+IqJ
5SQHAPlMXXxvxk8a6lD804AHGzuIilC93eg7F4Mt3R4veuFDVrtLlwUptoCl+JmwNFvAvNqmZiN8
c3qoj0zaVny/CpnYNZb5muzhK69LWo/TLs7X4MVNlMXWPxIUpyTJzqYSYQrOFkuQ3NhnXMiSVN4k
5/GRAxhVIPVgtU89FQZ+zVV7SG58g2q7usDqumzteJD9BYbXahRJZ7WVGOQoufentd/dHQiLIJhb
9shNcMGJIxbtcvcUZUf1ysSGWgrfmqk0thlnoB8OPZ8Hx7gbZn5WeDWsqcU/rV2LJidZSYsFisbm
NH/Y2QeuJeTmUuUuRXVPaUkH8ria8ULnuK3JR+gkAstDyHvIW9GnntTZQQMgs87PnXw/NhyARL9S
As3nj5XJvtyMGgLYY38PwPCMCqXbWxDz6yPmyvvEZBrBxoimVxu7m/xOhy2bE+MNUY1zU5FTu52v
FvqZSLIa/mj/5r5JEd1lipHg2fcOM04Cyw9fUXHy5Uz2tkqV7USc3D5p1yEmF7r7/pmcX/4hqIX8
CbZZulxUyGFAM/FUJDUx1gTfsTyumdZ+QeYCecc47hQXD7aLXr0yZ7zo8UQLauBAHyhfQN5I69Vx
MLm4ChEvBNsQTF/WX0+4Uvl7BQ1oS7NM//yWR+uPKTiJsORvCBuuRpOYXFFdsWAeHQKeHiJsmUhb
MvcDlid/3O8bPy265OFeMXR6pVJhCZWROVegqOUxIzRn8E4AYeUCH4k0u1uwR9fS0BaNL9WkPCQx
Bz4tpc8IMUOVyqJeYlcvIo/R/jHm77a+HiS0ico7uESJSFwu7RUXQLZJDod3YTauf/fmiwjKkl9B
/VcZz21/fhQaUIoqsiI4W/tP7zw+E2CtGb0AMBZ9MhueaKKzX5pm80G4bmfBqNRl/Bt0GZk6x1Ob
QNMbpzI7y7xa3ykcz7NTeqelvm4Syv3S5Lc+y4PVgigx9snql1UJXEgXRbv3TS7cmOwW3hxxZY48
6QkufYikAze6oiF2+8A0C7C9Zauijd3JVauZJsnumJnFh1sQIPnJKy7S3BwtufzpucO1YcYtYYIq
1OqN0uUmQvE0l4swk37zENN6/yGFj3YrjufJFIs1xSfb/zvPG3UHxQBBl5OeN7/2Fshk1yjquB35
UeIeXVvu65F1EZYdieENUsXK7oFiMIzVlbB2IWfXsc63L0BO4gzPIm3TgilBiXNJUDHKHDPExrsE
8Sm3Ftz9FYN6hWynKwo7hNQDRF9X8SnvUwh3CRxIU3xjXoNexOTf8jXYZ1UXAcLVJzgQzdQnQBEa
Ct/J1JdjzOb4rlrc0MetPm7BVR2xRY3QXv5SUyYHBvkne7pJif5bt2GsoiRhsc+6xxq4/DTuLWIE
2t95VDfLGCWmc2bHUtZE3n/xiVWnvmorSzMOQC1ElveYMfH2qFrx+aS//9KKupdPcb1MFVoW8xVG
sKBzUd/0E+PCNfu//eQCkxFbwz/fRhEOG0im9+mMV+JXeeqVd/7idY5ZdKAgU/tDglhKKonJNi41
QHwbgkgzJ8nOsF6k6xYnkYFwUco6inyN8LIsEenM99bphBHvA/F7JX1zjnlbOCBGjws5VmHQPgUI
/Esdks4EugnyJAuvPZd88AGz0OO2XyuO4UeUmKO1O8LPhupC9raUhyI1clHUACC232ATDWfpsM7q
FFiW1gxH6h8dC6qFLvJIZE9QOX9PjaTi17PGXRrLYT1+zvUEd83dzZAMBs0ympslETSMYyFID/9Y
uRipqA8wDEJjCFBbSTI09RYo5ZK+2J1NqmHrQ8HdPSXGt9rI9YxTGm/ngTEne+e6zNN2CugvZGPs
8uST7oQOE4601kdJt2C/UnycwXZN+dakuaEMq0phxGTb8q6l6dU1nWwOR8XulFqUUlYDDEyoztUd
2VtYJLqQJ5AnSH0aTgvDI/R4CnRrcgHyJRjIMdkuxSGyZKZeargI1ikcUNMzrmDfvcCyKZaWxrTk
eoC7cr0DE8VjRnOj8VyTTXFlmXf0X3fozl216ADewDopqi429rtZD8fCYtrvUkZE4RS9/uEHJlZe
q2pab9pfoGVKOoRJnTSUVg1IOxTS3P7kVXx8tO93CHF+8TwMiKWN23wR6lVMFTnTvWjNmpWNGSEs
4pdjwDE9jrmoe/YW1gumluWq//a40svfowkD5nBnC2WHdiaOmlU9e/j9c+lPlpsiwE9szcB+TLKc
JC72iSV40kh2HMWPm9aEVN8hEacrAtQ6z3VcVu1biP3ndUAv1X6g+hKS+UVlsjdG1tDcBCzoSFcB
O/mFGvcfF27xT0SE9NSXgUJJrIc15X0C0kA5QPVD6ZjPimQnMsuOYhZV/ShJYO0W4cbDSvhbrYj4
ISGIz/8olCnnueuXKdOfaABAj5HL7hGAUEurD4uAHGW8eaT4CxSH7tu+7Vjqv4EcMgyV2qfQ/HSg
yUiZoSjeEuqZHX1FKy3HjP0uww0m0f9LQYYa/7HcMfQzJ4bnM3JVbEk75omyYbYM02MHPhWS5m3w
NYSpa5bNJttF8F0rkTFzDIfmjB5ojHSa1sdGQEjSPDpVhTKHmzaAW6n5Wf+1x8upRIsLvpbOGdJY
S7GvOu433kqs1I3hWjk4iJsDIw147AxsrlQAbfOISViRb15c0eTanWdbijVfHLxvqIzNkRgA7gRh
8QFyCVyiLmmkAa10qaBXefeRchkBDqPFUWMj41fIVGtYkERug2Ufe3tKnFB8ypx9/uyKdeZPeN8M
Nkry/Q+susgPIBL3+7OMK2CdQNT3eiqWJRdUkc6RQRsvbfTtcALWQXYLBrDtNPXP25MkbXkRxHDI
C8ihzYSt5oaEcYO7+43LQ4NEJWBeLE5qbG61xS36kGQUdyjlXbllJstHzCPXJX08RnZSgFvlST+A
H4HWq3trUDb40mvELXTawXPw8mi33TJwwUpp+9+64beHGUFyhCHObc/W55Ie8IdFshdCSSgSuqZn
8JgMQ9NnS5xGYZqQ6FWoIAflCNREYFyqW4KZmJOhWsWlQOPJRANIMkv/bHaENMjg+mrmvXLAgGeD
yVnfxgXd3euxuT/dHHt064kZ8+gvp4zy7ZehV+dYrRXZm0lsudlrtLyHe1Rr0zVeK8bywTBHoNE4
VpYpzZNhMWXOxOfVgOC1L29JoAe9nHAIDD4iFas/ppAqtxVpZr9S9kyaio1ojvhsTF7oxFC1ZX+8
b8zdgfFw9pPKRtINRyFWTduFJmC1I8Ew7wLU071Xa2r0gApbkXfLeocMQ5upGTLiEFxbNd/JPcR/
cJk+ZXSoxe9GgHsy8/ggFv9YxStiMyCci+ToDnKrH8q+5pSYdDq78CkkkNL/sXTbKAC4izmN/YEU
qhMN7n480AYfFanpDuKSaVY5Q84JQ40SfMf0wz4zs3ET2Qc+Ouyj06KS6vGkaNK4k6yNM6s4fARu
f1gyX2d4lLFee4oOVrLbDcJE1uqUNxEJMdiJzkXZT1xXcuH2TA0TL/a8AKKhKFfTX5pPlaQixrc7
BfendjorKp1U2fkLj2GVC9MAbaNDMpH+PZLx4mCz6qIX2Qvw8Zg6B7x60GOVOeFb8nR46+DJkJwE
hOvQeqz3/rjdpTTiMO8ETcH5pPC1lDrR3MROWMLH8mwbHS17M0F40uvzcaDKZ6MKHDOo+k5oyH5n
ISn+qX545+xvU2xavWxO196tyHTHaOEXe7BWtcyNlh2vyarb9tdIVJKBN0gShAhnGwurwMS5Ke5y
G0rUX0XuWmegKmH6qGlappWyInnn2xQm4yrlKBIoCkDZuGTPLQTTbdbuPkUm0Evhy3Uwz5/VGQ1z
PRhOuMT2YFiuAN0s5ZPftF1A+/j0rOWwg06UCZaiZq/i405MYKKr5hkehxJyWucozYTWGI3ydgPO
cmKEfg9cFJX2JfbQNU9nWotQRw2eVuWT9TkGU9lo7YJ56+k4a//XI4Jj6hFfr9kMMJLH8LhRyTDD
nm1+z1AH+DAKTMUvLkw/iOdhxsU3cku90vgBshKHcI+cgdiocarvqxRCW46UHhfJRgVbrhQAVzHd
0xmHn+wubZlMxNug25k1HjULmUXwCY4lMfn8B4Q85E+e1domuIhnHyZ/R0u9NBwR4MoclcDMdW8t
B7tJeMjaAnMaBCDgKvxBo6f55CkiySMq1KKE+iOAmXVVaBS3YjNHoV0IM3iR1kpxiNg3VW8DZ/TL
99EK5/k0bPQV/l6M/dBINg+0o666l4/VPJdj2pV1VyeYZlmvXKJiS7QdnK3c9+0OAfhzoSFa9ou/
ZDWbv/aaQ1YY6mEb+y8426Bqyl0nuXI50zKn1LvCN0veKbtoMCKZ3O8KdBS+4J1WbdW2vuqnrFHj
rdKLaH9TbdZrGglPEjdS68pLLzov7Ox41SWeWJ2dsCxjcb2DHXBhA3aEoBzVqqcpQkaJY7XrSyE6
AaKPEgIxVM5ozw6Zdq3vifZVP/tZ7IwrB6BSW0rtktZlU/4ypXm8Cp3u+t9hOZcEdVo32/DaLXp2
GESgXoRubmRgb/7zUW3E4qXLZlPPiWWkp4HGDQjw+DJl/emXPJirokkzWoct0LH8QYp6LiFbF9Nd
ERTYpiuu/v6c2O6GWwM2BE4UwHurn0b4d19Wdg/nTWmwMtdc65C7Hw16UuICrN8cxBsLvxlsh1TK
1fCBUvFzbveJ10vLTYpEx3jFnjoxIoqgNQa8TwW5BE6OIQgKISTwp1+TtpqFjQXycLOqGTCKJEjK
0UT8a2/Q/J4NJQjzHMxtWn0pLIHwjNtpxlOdPPtenQI+rmxFS+DCqh/RAEaxvrOtjGranrhUntgu
zYQFo3p7ov5xqAa5WjKNVXvZRS1SmrpfMinCi3sgtNTK7ZnFSLIbnf0sDcfvs5bQgF4tiWXYEm4m
gH3pvopfedi1gNLGcJNGgFXnfAHVhinOxVcBG6M6x99mZZMKBfNhrDR5FVV4UBXKgcS2pglDITMP
hgMit7uutj192op3n1QpVQ+FpxOvnM+d4jwcO3ZUJ6KWuyS1vJKN/KSYYvRj+wu7R9luQlui4JNJ
pkkL3qCcNO7C0Hs9l9rhfsurfUQyYOcbFVTpggFtDE4fOqJ6nlRJHsaHNHL4yNb7G4ORHcy4Du8U
uXvqBqhicsITnfPhtAFfnUEZcXGH29o/Vl4Y7szrczhY8hAXW6m7ENF3IosUK4JXHvTE7Db5VCPh
xVhc2EOOyQKL+VdDGh/e381vNoHv1cMEcF6Br8wnn3TgGIOeuV/xdfVKsugB3xSTNyq0nw666nIx
Sbwu+jdZReYqpFmRoGsz5jhXFIO8eYMOQUC7DGXRfD6WSW2Jwd9C+Ib5czCUr6slDkxRuOdaeyYv
Pg6Dk8L8qoCt3e9o5M+9cqQFAb+OsBrj92APs7tCi5TQmUHZ348r3JtPBRh0Uon0aXC0qiD8ZtZj
8UST2+/yqEdg7zoFdJR6aQmhR5h4f08payvRW3QkVzbuS/o0hAq/O9btsAWMCSnEXpMlAHXiF1WQ
iCS2GTd7fgAjzH8XkpAo4jf+CS4MtIwrzWqqL2xF/DazULTXN64WsI6Vz+FV2QCxVRHn2HG3RSF7
lVnV5tcjpSsVIWl7nwX3V/IIfmEpVSQNOLW5Pc0lvUHVbqrJbQUV/RlpNTOs4ZhTrPC4lJzw5U93
Dik+xt1UP4LXMZdDjOI2QNp9q+RRqcFRUKZpYyIHSp784tVrv+FIYkn9ob96lOiFETIHaeMrZogp
b+TdJSxrIAUoTX+qXSfnG4ED8X3pgib44AlwIVYgruv4/GPx0uXPreDHVzkA4opY1s4nLKm8t/cE
ch6Tj+1WyY3mfBFngbj/RjXM+z+PHV7s2OlbOizkhAK0tDYu2O3L44iIit/KGgu3NoqVHfWkNZub
pY1PWAKRV+1yQyHAyflxsO7eVGUrHyEju+gNVpOfOC/tCoH3j8W9H8krAF8/cBU2jiZWDW54eveM
lKpSNBPb6Ttd/ZJENDgyrlkTOrQuE168yUgHYi2+QAuJ85GYgKxuSvaHcQc89HsNVXu6SMjtV/6d
PXxPkhWHwUA7jV/9ME9l/V1NN+a2k7eAg18o6frWHH2aEQi+aonCPbeBtYlEnQcm1ANqo5oY1HNv
Sgb7Vqu4TRm/7gU/Ercg5gRKca7kkx5wjfz0qbvaPmKxdedJ4o6gOt5tTbvEKGNfqlK+cpf9Hryo
ShWwbJtSjfZBYHwcZcPK5i0YHiuW5/fZQP6ONzfnZ6ms475H6fupoaczF2mDWqHz9b7ByT/mCbaE
dqHdyv2tj9WL5+r4xYgsrv2jXd2W8gSkMHWX5nOcG1ahqSoFVd3aWBZqBnVX1yf4lytlduepR3nG
aeNed0adjTJUOzz1yVHpaeAIFb/sdMmOg6aY+jBkwb2uI13OF85W6x6wEq75D2dozCsfY7I2WlUw
/iXO/QpEmron0AzmKVq/MSUnTSFy1dHEvv5SBzWzZEO7lvfelcANkxMWkf+Uts44Vh0QHsMwUwq5
jgtfr6NeR2YFq6ryeK1EFlLQut4rA+/+PFaLqMG/WFrbs/3N9pnIcFSV2wmERsd3zt9NsYsxp2Xr
9ExkfBgA09MWl3Z2wkX+mpXmjy0gG+YBu17lVF7olnVZNHGlZ4S4qHpNMpwNTmZCo4LmcEKNyZxB
rchLVkNs4JDl1e45/InekqusTN1w+JKX6xtXkbLo7BAUObpUCAo6BXXqiig10k5M8DwdEHS9RLPD
vax+Gkl14NloeEzB3Uz8wx6W+Hl2fsgy4k2fx8UmEnn+0E5le0JfopZGHzv4iS11pF5UG/M53gBB
JTfbDgD8/WGT4/sujrH8e+5+lnQql8fV7ZwsoTyNiD84nsFOObtLzFeH5JIpe0qBMU5LiC7m+E9o
m0NyK5msrvj2AlyK1dtoWrAXFrozQ3oGUkk00z2W8Y2+Pm2bEFw5t+ipVyeHaHE+ESWqfDJKQVI+
jFxce4K9dHuNWgsdpPfW4J+h47pXurGePV9YH+MhGQUPB5/XDzw/7Uy56I8kat4hpxm4S7rMHKlB
28Qvpzrw0Pq8ZNjAyVszjpuwVQzcUOpFMuxAj7rzqX1coMPaRP8T90Ohe+k7eW9CisSGQ6D1rsCc
a6xHrJqocdgz8IOgPicKBpHyt6VPhUOB94NB7D//jS6zmF7zUiK5WedbhT+imS5xpVXBlOJm7AtH
pEEZVkUa0TSHtQB7RQCRkeltRHhZ3UJSHOaR87y+aAT1+0cLCAhqwLKKuOyFR/3HIvX/S9Z0VpN1
rRzAuaz9CZp2qFDpib8YRM8H4imwo9RcPGOH9MP5rQrGximVSc/af1GmW62PHlTQxP7MK2z/CIK/
73Vr726eNin40BOa7ajU9cQPtDyJTx3PdAi9oIrFfb2FCsYFRRaTqciqOfFojX28GoIldfHiQpwG
oP2R0X9K2XB7O+dBa1ezd11oiFpWBdv7boSNzbwCGbikUO6CmLMPyuQtqGk51ilpquFfWTccAa+h
6wtrPgaMi1DFubFcAMToSHVwIwiTx0a6wKvVCusj7ZtkiDJT6g3y6l9t2L5ZBuPII8+aCiDmuqNd
rkFFm5D2yHhQWJC4btUfQVte6fw3coGR32ec5Y6+WFjaxRcLb6M50kxKjsNYunFoLb70ZmCWIPad
g/bCm9I1aYF/wwUfO8JVEz1ATzZz7CrvVO0hUvkg+nIwSCfshDYOneP0OrLqSCYij+WbgYyjEEi9
WxIbOkOYPe3WirLG6F1e6FtKx7NgI236gYD9GVidAy1CIZH8rZ1DeO9WYf+yV3vPRtZujATUgehO
oNklXwMPl9Lsf3SiwlnhEPcuFZe6HnHVUpveSCeIjb+7rdWNhHTRsbjcj5WIQXYgeZ19epLOE1lH
OGFdnhekYqJOdNv1lD0qeD5BlchJIORXFyu36MJtuxXnaRDXT9ZXs9TNQD/HFrDcsWQGhmG4UhG5
FE1+KrbCX7tyMuf8P7PrNsSXncQmRzRqGm78DpAvdIPkP76H5m/H8xLXtjXIEm0LX5gJgolyND1A
/Jh51AHfjBtr3a0M2cFQAbqtS3Jdp7M74+lcJ4FsMkvwPMKbho4wcabk6mkE2nUzeIIIh3WKi7qr
b+MHLOMdBvRO9LvuBEEUrqO84fQv2EjZf965ahZENznYvfqFkrIbvBhrekwv0Q/JAJJ57rRbLVF9
NhU6VVhLX7BKsxJKq80Dhi1JYt0ae9o8uN8pgXJg/JeFjTgCoEtUecwrpIyNYJdlo2S4hFThyA+B
D1vMxbKBAiP22iRcFkmLeT7E65oeO3lVo0OzD6VH8xkOw+Y3j/fNDdZqQMUvTycsmbMfOrQhFUDD
E13EXAupWAA7H1l4LvNFHuC8DhShoAJk0vN13gPlM3YhObIQytSfHWi+pw0O9uK00p8S4Y4FKQCi
iFDHjVjpl2TI7qoEfLx2QSkc85170iaysDD9Z5I24ab2fpFeAElFtH8bmcmci4PNc7xXuCVJy2N2
NdweTuX4sqJrtiUhs3OC3sfPtG0iCCjeWIBG0XdU7c0w0C5jcl5fIEqyGq/H31W3mSNxpNSFya6b
0VD+m64Ims0TBxzN5ivYLZaYwWf5FdMaHdsvbpKH1hc4rmeF9QaTcxVFdRh64MA2c1PCf3zQ4GmS
qkqWldalzOgRQUY7otaK/YSeb5/bejFVmqV8h3gTI1i8Vxo/rivvyM841kWSO9+3arXYZQpWgCya
V3noG+wBRlbEsHax8u8MVTHZdi+sGkp8y6ot/7yyYND8II8oQBy31ylKJeu9t2eVBfzo3kzhUlNb
ly0TlCNcbnkc6CvT0IFODKtRIh9U9g6nrxCJm71/SexQuuOL2uZntpYbkhWxLGJFK+ysfzF9Ap+q
XaM7MLfELohkU5CPKS7jXMA1e45rXoVC0B341W2dyuIEIC5Nnynw555uw2iDDmnn9SCi0RthHlS8
WrLz5zjPUtB8OLw+3246avwyl3Bwk3uylxrJ0k9plmxtkVF98ntZfaLrMpwrER6Mbd8rZP/Z36UN
644PRSZXtw3GwW0DIX5TxqOJYgKFqy4VW/Vb3Rq+Uy0nByz6lOgN+65jPjR0joGRoNJ+ghgNbjk/
g+1h2IvZvJQW/utG03omB9qhfrSSTTV1uI70iN0sABnY8qG+AXz8HEDKy2hctCxVa2yegU6xaMSh
YBQksAP2FpFZsmUyHDDKJH/tcpnMUjp+tbqbH8phUFX/QpAzq/TNz1IXpAM4xQ+duJc/Bmj/mo8O
+fhC/ksqQ2UN5kERlbrVRZshnFyQjx+NR70weC+mH2NN2QaqOs5LeTuJZZ4y0i43H5sx7KjpkOIv
lDXpeGAlAzn9T0kAKNBRyAp9VIgcqR50i+Q2YhGJ8VzMA2p3senOmek4yBhDlY/TZ+n+kpczSeaB
nSxxHIvGvn+0DqKOj4cfHHbm7sEpUgw4UlcnunZjAJ7hZtLTc8rAbXm156RF3IL3K+3FevFrzM2Y
gyrD+Um8289g/sh+qY8MuR9zWB/+34sogE2Lwwx7ykR+Lt1UtIGgd+FxHVa/TvvfWl9Ssl0GI4RG
wZbOujMhFPUaVbOfpFyit0kNJokfZsEFWs9M9/GIEKGMMAqKeVmy+Gf8PkDIsnR63tp/HKVUeFGb
PIUo1ShkYgUr00BZ5jCjoOHwrludk2Dhx095pCw2HeXpST/4w3VX8IrYYvjVzLKSamzWDxbilJWJ
cV0IxVPcK5cS8Dubvx7TbpSurK6mQNFOG5lBHLqVUU2A0AChlMQOoXEWgczwSuIKaJx3ugOqR8qx
puUQKQgl4dc5Jchm4lPyNTYBAA7SEfPKsm+Qma/t75cgnpFoSMHMiM0dAm3q4BWTalwaXgEoNqGv
/OX1UwB27R/DcS1F7/5gdz6dU+devUewKa5vBT1lY7nC/l3vjJCNoWVFxwX8IqFYhri6diH0NGdt
rPpCmLAkDZulvbOh7Nz9SoVuR2Ig5nFTI7KCXmtmegLPB32UVZ/lD0g9kBVuwXv+oGa/YksZCb7s
R4Itu0n++zmsG4910/Tdc07M2QxUeD1G6BVBqYcB+vGUYQwKhmAatjXB9XJgR0HZhy4pJoeUDccX
8h3YmAtCmJ0JKBTxtrrECjW4KWb65ty2W4Nuo/DG28otXpdSr6WfSnx5dK7lL1P1TsWHLrh+c/GO
uPGivEhL3zgDnUwd/FPiUwkuRTFbA1JvBtTsRNqOAIqS7rqmpJhRqlar4lHTeiFpqAfjhBsfg2yg
XnG/+jow4H813n1TMy45o5g3df9aqAr3Q5VMXFEPquILzCgqLiB0QOoo5qku7F8y+Z8sKxaWNrOa
NJpy9JJVWfpu+TruvKP+SkpdlFTVjVRQt5y+apem8oLjbemQI1y0vtH5Pl05x5QQlC9+2+JKvYGL
UUVCaY1raiJbU5mq/MwnzIt8NBDH+zTvKrOaDuzJLlSKAgUUV2zU4VSULT4GcnsaoQawW/b+OVoN
mV/e8zo5MZcUAj85vPxdHH8yBpeINz+Azx3oCbyQDLvrQO8JGaJjRXWBASB3/oyqifLIj29/HR+Y
d/luT0GY7dYD7Qow4T2Q/A0gEs/ruzS0h1W97FOTmThKNlIjtg73kRKO6DvEBaat4yaiscnz/6cG
ab8kKveu48py1xnkAO7RxmarertkaPHefToQoeHqySHdwbAWEhCiaxp8NxbVZcxiSy/TIVy8XkSe
Q8jHFeHqwwmhfA7wi2sh0g8CKHzW1y8vDdDQq9x8yNM22qCQ10Q/j/STEwnUkebtI++mo/kpuD1T
q0fidhyjB+U2n8jqOvirZQ37KbApwAqXpb8EEXn3s4NvKSFq4FlO7GQCDTkIlUOWSTFtBbAaYn3V
Kyj9remcL3XU/0FHIAaDmUBuIV3jUzn8OL7/YSjV+37GHsxaVWwbTIQGwUDdRZpGL4VSCWlZuPYD
8W7chTTdRgw/wA4qqPQ8iZsD1FIIcyBh1DkoBq6cZFjCrO2UdX2oijwiqsHOMJWtvnCebK35OhGz
jCo8cFjX3V3H46l6wVqvBfTcVedX5Ywiipu2CXBGdGofWYydQcCABiSQtXWMfc+6tsPy74qYOti4
LJFMA9EEwoCme1yCTj9Rb2FhTqS7Uq9RE3zqmgsWec1HSpFLwtzSRLAOxqyx+SA8EJvRjZ33YvII
WPjEwXHEz6FaERaWXz6B7Na3ySZ14YakOAtd6PHzZvIMcZ1XpvezL1yFu8gR1ovdBfC0taMDKMoD
eq3oJqjudHCIJuzPJhqwvzYUEUHF2y7aRU/DUZNiDmZQgysEMlLKOmpgmEnfb0PVmp3sYNHKzUrV
Zo8+vZhMrX2eBmOV1yPeDjfQAevG+gvn+OgssizV+n+KjQ9UyTTrEh7SNLH2OThYtPKadBZwIMkc
MOrXC1DvtOnIaYKAbX6GEKN0nA83h+pLWyxR3QoJWria3N+0A/feudXUC9BHybwK0sE5EEVElHkE
1XSVuawQOrP5chmq0FVyFNoU3cVnLi0LoP0ozk7Hy3FrmOSsFnUYWBZkX3p+2YpeMTUdB/ezRexe
tp3dBKTehX28X96VXy0hlppayln4caNz06eHpl0N40hCp7PB7TpdRp2/I79p/sL9rDjDyrUim8Y7
lJORGDEjao2HzM1RD+dg1iJ9+EFxQh6++P+Fb5jOWhLP0UAb89My+OhgiCTf/lA9Ow7FO+a96NL3
5X7VHuS2vfUEP1d8avEs6DJKC4AqjdjNqSvUFVh9PFMOGAzopQfS8WzYYr6vks7JHDb2mKJGuWFN
gmxGY75R0rAjlET6XIdG3JGhrB5mZyYILT/PuOBAKjrxmTDGKsrhjmpv2mtjln7ueOjUELHtjt+m
XYkeI1/VV6Qm8vasq7Xj6oy8HFbpWowinPKivsVxT8ll9agJxafw8DymgthjilrD1ONBdZi8Ks+z
5dXXslkhjBrhGujvP5t4oBi5P6QdntuicGNUbbaYMtT3iq7sig2I6ctn+FZDat7ppgcgoNe973Zf
APR2UgS0rBsbgV8U3ICJP1cIqU5QGrh+PSZQlEBeayYfjmFiWuQTqm4z3RW6WEZ9moD97iA4iMLh
0HP+NKQgZ/aXn57noLYkjmGfzR/zO4kSXryNkYoS6TYwxw3LFmmw2yi8x2zh/pXeEHT4tFSNMS71
6woxjiR805KrqeO8H3dmKIVVT76pAmmDeWWiy9xgyJNznSzn/lVMq7NALVopwCDe7Hy55YipBJTr
rtZNcqVnkq/FgKkTMjHcWkqtQNHaKbOuGVzRwK8tFjB8IvVDp53dKlk//Bu5UBpQBEK7M8fbRtAu
Q070VxJOBQdLmQAxBk5yaH4cKiVfA+opqj8UJmYtJGHW0fXJMNGQrSt7p90lpIYYmqDazABo9h6h
+PPysLgM/eQtvAjLV/KN89yqVaRY9bM3tyEiKCGy/7RKcETaPytIzk3o16Mx7RXYdoNviO/GUNl0
YOzuSJKd3wuvEinEbjvJriKSji0eREJQIcTDFBCrLC4DCB4ZSJmKTZpLlT3lVj28dmZxkKOvtrgL
nYptW1Z0b3gvmdPXRSPYcMhqI314A6ZyV3Je5uWHSrXAsNia/IPeWYJR0LWfuXxkR3Hxi2LjEh2v
t1EFjfLjH+22yU0pz0fTYpiWyIwzYClhwRUfTX6G4EcYeV5wIXXdPA6hnAJhoa4uG4N9QJYwQ72h
LGRJuvEb1J+sVIsDXZypgPiuduTHxDgFsXINeK2/6g+ab2h76StRNgF8evy+/GFM5cFqBp0RzX77
wOxTVqCJBt7C2T8iXs8j5DHHG4+eIBf18Fw5rIHJN7nXUTPpvSFUVgXGSPc1tUr82Yzq1u34Vnye
R5QK64CuBtgbdEMHA+yvH3wRgd5N8354YLJa7tA1XxuFdr/D75AJs7BGUpU1irD7rtbbAWQ37fwc
MwxKr9A6WztY4Pkr/ZGn8OGKRrGrW9F5TKYucWyEOQ89qSutlfYOdsAb5AWZDBtmWbgbbK+FhVdi
1YktOlbSBk4w6tdQ/XAijAWL/luQFyOCX4PvaQtaPOB5gHerbc4aUo2w0L0jLxKGqM/b/k+B6+Uq
fJ3qnpelxigLQgNZZ0cALtjau/TATXQkR6/XT6RxKXT4BgNv2FYTtQN1rDoj6yB2NgrHhs7IEBJ6
y4czDzVpiyq1inWoSBvu0eBgJmZVnIyH47RsC+6PrwnTQce55pD6QDH5t30XCOpHZEypkIHyrh80
URrvmkJcGrbjARxRCyTGPl+8EiEcp9aHHgDzdP/6BYSs+EMIscp5HGE/jzshBIBBmJ4PrrnHIjL8
xBg8POmq16H5vY7A2PUD0JxZqArVJ3t8ev2Ib1z56Yq34FOi3qhi4kgbTLNIN8IrhTCZXwU3Cbru
ngnKzR9dJc53F3R9V1L0Z9o/BVX1vZZ0mAuAy4e3ntGWW4EAN6M4K7MHJFmTpfiKqdtM78UI5NUD
8MAQUjCJeVjsnYXW5YpQMZd0HEMkgWWP9hKOwDjZKfDIkz09F995Dj5rmBzuXHCZkwRyBI/1hJvB
JCZB0z0zGiKNoetn/+aExKZtH/TtOjrNlhoDgFvXFMhEhkIvO0AceuiO32RDbMsJ0jrt+fCmlNEg
45wiAp6IvqaqEnkWHhSA0HiSgsZYHafyhMwN2A6Taj4HnQ8IUyC4ZYF2wjFejS+JCG/xRh+coGJ4
JQBLuado7Rqo/8LXZ0qGdfEzkPDc5SE1mqYfaMQD0V4VGSYjei+74M/mCTYcyJ4GmraRqBPzR4l/
2CDmemVfPuU2hf5S0K+yafC52R3X+ihcQKnnx0yMa/PXz7dJIPiDVMiLevSz/g2UyeORUYXSaOKQ
YimovAn07lQM0icX8q19hxQfbEsoRm1Q9HiTQIXC/4i2hra1eEvEx0fAESIwwe0TR0yJp3NDgg9k
W71giUHe7uQawgW5O6ufwTgk92iS4ZF6Lzzv8WxUY6FCxjFsr9wMFi/uFSH6JSMKGpK8vMI8tGmQ
Dd/327r11yq2pb8YB9dpJ4B8O2em3SoX8//ocA0+9txH1NAxVC6+CffmY1N/IqrlRWfMcoyYMeVa
t0GrgQv+eBLboDFhO0fmE0eFxWQKLwY7ERrRGxR521UZQV6Hk6jwDCZX/TxD44BGIgTNkFHnInDW
rHXPKQ8njwBcJqyPlQvOcmkuRy+kpg4spZaXtIvxD8wZvTSSpRfCuUevKkbD4jp/DxlbNH0OYXGu
pBTmgFZW8vYpaGTP8LEZXbqJW3TfIbUEnDmhz8ZHrIqRl6DachAq+bpzowy4J4XgqzBA/cHGp0MG
lBRtzZavhC3TVD3c41IcBvN7RbPtbnumqNg1bYpHX5+Pp600StH+J3+JUKbJfz9zvk5qNIwxye+Q
MTearMUqLl5K/SjkcmC3Jsi65CBJN3pd5AJGhMesNBdyHoNx0Z+BS1Zn+ay5KG0etwbN06FaQswv
QkbtGMZByKCVrvZgvGlGmyLxO8G25liPcT/ZEYicylIArTKqS5OWph3/6an64SXowFd1Fbh40OO5
hqJPcurAgkJuBfRbEP1Yuab+WHKZfM3Qqhs01oS7N2hooW0TCvyzmG9OrMsr8L46P1/nMWLqQvl8
F8FNKOW/HyEbgTU6KFAMYoT2oqXUK5iFs8zWZud35dEN19dqYHb9TGwbInNET0yG193jsySeKdw2
IxOUHsy2Fj5jSUxHKddmOfWYre/c2AlhHGpqYFyV9tfyPIQxlWDV0JNruLIkAq31Zc68LpyuvFHz
6zY38T+f3teJJ3BozjOAwrGtaZKWAKTypuZlET/Q8gd9FhuSL+7kHeZNUl8VG62XYd9fJYpXh8jK
zC0D1wbedBrpwSpNqCcNAH0wgQJNiBmuV5NqSGXWtDv/pTr2TgZR2Bv/5+hawMrCI0ob7ohOMMyG
bDgmPZjPmStM3P25VhCeWen3zM50HRZBkePClprX+dGSyD3iHHTvwZIFLPmImtexsoBjsKaaQBXU
2JTP2/XCakVEF0w0U6qLVfRSVi6DmUQHh0/AquleV4GYpJBkXSwo7SKfJD263GnlegMSusscTLE1
aighCuG9HREznLGbd1hF6GEH0qcqWHsKD9iqL94R2r9PS8/gnUh1QA6gV9FMoPIEwGOVpG3plE/b
W4hVOsoxlS+ANmndtF7fr3mGCo9tSAyUzXnSn5pSbgcoXu8UJQbxDko/OEK/7DNgDEMQCgbdxTxn
UKgYr6qt3bDIoG24soedzDmonrdEqQbUOUcXZxUa/i/Ool52+sgmK50DZtfuelQiFiCkZgTkdU/N
ni6g89bbzGQA65RHrKMnzHAaL/V3h8SQTXIft80ZrrKz8gaC8TYj0TA9VuVHVuv6jWTq8MeOc02H
9dHMRWHsUF4p2Y189kStZmj7y3J5PRMaBatc8fyk8l/yW474h65Fate8thculaJgmNuO5ajHOUDN
Hu0tzk1pPOHCVeBlaXG68uqx1px1NhUDR43d6orufIDDPoh44lKh6A9/fJm4DzJqTjaVgNcGV2d2
PJvGgusTfzLWyLBa0c+lsu/umnnSu6TY1um9sZaVBelP4GPKQRNJqWDf4kqg9wsTo5Udb4aGH8gl
QsKDzI6j8j7BwD6f0KPY6VcLNrQNvxmoJHaUySZraf64fM2tBmjsaC8D4ljGSgfqUfop4GMlfWXy
UvSM4t9iH0Clqt2NFPoDj9cxQCBlUgHwBAgUCMNXPlgRLYkXXu9Kn/aERgG8qAFjHQWxosmBa5gL
WnUv4twMCvBIbDZXmROdDX6F73XpnfXC4D3ZEoDcJL28OSSKE1uA42m3vkRQDjcefayq1YBCEisv
/9l9ImhYqvDTOjM9leo2r6uBm2BMfZwGsYcRQAvLM0rSDmbBR65SbsDSzXTJ/Fr44AUW5MAy+FS8
EBpaUyun7Tf/TlTmswhXmdkRRB2i/uXX8ftwKUKeQ9Q1JnQsXzfPHpqKBlmpZ2B5xHY9NjhvkrHk
BlSnp1jPJQlYqNbdhpJ9043p/1tq0iY9E97aZeNYun9l56y9whAdoK/Gd0hAw+hiKPLNwIeMlGoC
GFYHlRVX6RgxXiBGq6919d25kka+1qf7mhsS5eZHeMvx+CiAX5Ipp2TR8vL6DEmMTI4JmNGE3jBd
NxzSAdzRuj3oFOmYQ3mlm+z9x220uk3L83iC8m2syiCVR1RGJEvbS/ruvXB7BjGqAv4zJhBWs+4d
CWkHfX5Moe5W+HgqqQTUJJLe4BMQ3/uoEa2pgiM8fYiq/pwgQyb1nie22n0eYaZvNwhFdZSXpn5W
BZ0d4k99wIBLIpHq4BNbz07qB36Jx9YpbWF2MSaUwl9ydSy4RXwuahadVNDq1Q7CjqBhnoW1ByJs
Y81wQDHs3UB1Sknagw58Pb3oDnf4Sjci3IRWgVTCpTkcOj349BL3K5zQ4HWpvNFxqAFsIy3jYXOP
5O0GG7KjNEAJtMs8i2EP1ziSStzIM+fGUpRm+y4oPkwf6vWostJLfSUO7G6YkDSg2u7/Dnf0aMAR
hhQ4RXv0drpJVKPa2CnOkP9XAbl301awRyODzmHOz+qbKqybFJ9fopv1TZbX2VieNED8Nu9ivTLT
6heYh+FNgb7xQkWMssZ+TqyTzDjmG/LVSZ/IAEyQUNiO9z4Fa1OdY/6+fnxefvAPSbl87V44CaxG
VoVUygH8k4aOCgQEho+4rzS3bqEyorsKTFFy9zxNJzWeDLx12qiSciUkqjUnSlTTEZeWo8uQhKbF
Y3KNYFSD28bx/Q/D4YILdZ6k7KMgDGP3zsD39Usx32E5GylAahcXHMYLHjdF09jKLj2nLhirm0Bs
CdnV6IVFOWfL0iQtcVunNk6fyrFxA8sa+OlZ4PAkd7oWB7EzKuaXQtWeFOVZrRS1jzSB6xC77w6P
XLXjcfXACIH4m/HE830Pkrrm0gW137Fn4hM6K1S4UURSz1D8fH0fHwnxgbEASHits2SITQiBVy0O
CUpojkggewiyBg9UiRL0rYZDNElc6APwd+k4mw5lIrQUkNgazGozI3dSi5WuqB6P1nYbQkB+yPaF
3Y9Wt65lIA90hx7yt+qU7Jc7+cw6ZtoZwVnGDKiysBnTwH8HXfZ2yjh8V8ne3P6OMc13kZGad8bG
PmAvZbKChdIUQJZmhN+Faj7YmKMnFg7iiX46GLsqeQt3r31Amqz63vQxvR9ISs6HYIxCW18VthVi
bzPXJ5gwwt5Czxf3km4Ea8QZ3mzzfyrXK/YcgYWHsqOEcajGv3bSCLok7ro7DsJKOfsXLEYYNPMz
Qt8lmnml3qzuRbFvzoGcVvyqgxLf2HuBdnZIsu156Qi4dfVqMX8Dm81eR2TRl/mL6fEfo+2w1ADQ
ZD56IiAaMVqH4x470fZhmEsBZ+n1YQfknzO8AuED9q9Fs3ylGzIImghWFu1pnyClVQgVycgGOhSf
500wq/DHXP3lEVDQGu1/bFc8bXLdHB9WHLU9U0XUxm2gWqcB5twifD804tqYDOh6F3m9lRGjB8mD
nbgUpQ/N+eYqazpwyscNQWPSHMBbF6ZG/6twuOPa9J9qYcClObT7TSbu5I6WtfqU/D60aBWDpSVV
2Gd5bxxNNgeRRnXl9BkPR/1bntka0mqPor+CReiqoCGTM6G9wZ/zzQnR5CliR1pSLZbWtUE1jlmO
tL0HNlH4P3XPp7JyEHWqGMup+r6FXnACI6thlmqgt/HaF/vVkGsUN4nlaBdEodPjdLenDDJcbV1Z
b9Gt9siSL1XTG+6g41FdGZ4tkq7j7qZCQsqz/LB/aotKzTpXmzRbxsI3BSJEDKOAY4bWtYKoSu9U
DoL//AoV+z/HAO2m5S67KcOIQsVXnhyEM0xct4Y6T0nIOXh4SH+yI4IxgkBQPjE27BHwIXeMMXSo
IjDcUoXDKA9sbtdzDGoGldaJfPM6f12ugIGMRJDdZMEaHxom+wcLtpRmtubWrx5riJvp2Tegk4Y+
4LmbLTwCuBwjdoczF8HKMPaIaN6W9GZVmrjXLqS1p9fdSvlVioFyqOetCbdB664A5jj8pJb6x91H
jA2e52TLIQk2N8uvQAmA5IqbFhVdCurF47Gqe4SNdFNHp3ZBnFd5HGiaQUmf8h/3yXwF9YQtHiru
JXv9Ggi0NSPNedbtZCLb6f4NvzDRMVAVqZMOyAUP2Iu7RYAFPgAKRsUiF0/XDTzXozVZJjFbs6SM
u4JjFfDUfmNBqbUdTgZiV5eBQPIEB2fsHSnp9/EycGehdJ+qPmEZn6CcSxJMvYFmz+PjAKYp9oJT
n3epCvDNgACejU2HFC5O1RiRTra0db7qHEb67LB6s4LRlChj2gYmpq6+L2JV4t3y3KSqA0Rfmw4P
LPOxcrR8WQUS5Q0gW0mQQvgujNqAH5PHun1CqZUHLwW8MywX3/G/uwvOG12DsWiXbqTywnM5QdBQ
7vK14+FfxAcu7kjroDvHTI4g3dG0daZFzWr5/gsUsUEJUve0aAxR8H/zgLBSNeQ0lgB4osiIULvQ
Tcf0fXVgci1vfyDpESN68OXUZSzvB3eo9cZsMc+aNh9GMN5YmJ9VANzQwjg4k2SXl9UgqwkgQCgs
TC60lqnBByBhIAsE3UhdIwTHDYcDU/qYB2c0TVKDgDnF9Ew+u/WhlroJEtYLoK56h2LmoMMALVMo
DxBntLquFWAKEGb4gH4+tTCRWhRLAOdg7TS89A68ZjHwSkA2BUHVA+3YnDVm0NrjgXE9/60JbfnC
gOBjAtmyoFEQUJ82824Zprw12tzIFp0YKb1tQ29RMLVrgmTcWU/0ScH/2buLVgLmmjbfAwkhAT9/
SDdoYbWl1tKmj6eWD/A0DkkA9aQh/x8P6dVOynkn3yxTOhQNHosgfgQMEnloR+tlDXIRrh+3L4BI
fDGF29sxZzn5n71a45t/2O4/ME7WXXt45pYOw0Sq9FDnGrQcedKX27iQBhOO5Y6rgZhoHexLm6Kw
mfzOIzCcysd2+dAOByZg20EftVUQkoyC8VG/JYTPZXbO5d2qdJ0FkxtYl7jiAVOtpQKUQ6yDmvoS
EMEofoaNk8h64SGOYG+jp/bJO3Egax6U0Ud+u5ylYETpKg06PKqJ88emlW+02xVbJncXzcDm0BXF
8cOqJS4+bMoBokOTSm/W3mdmM3nBQ0+tRceoGkIH/eTfOcImZdmoZILBb4sbkJjdz4gSEtyOZQwG
cM3uOEyofYqPmaAQdikikE7buVhWD7xFKGOvHpodr5r/3hWHJujDabm22S16kx+LQI/yCztL7elW
+vk1OBkw6/T61AUODoM5CP8wdhxDDQfjTgMJBF2T0RZQqkFg4Ga0YX1V/ApabbY9ZAMZAZQMiRQB
vl+SxPYi5YpdPPAauosZ6Pe49BkA7pZ3SQqZVte/VQ7//6YYkHt0TLY+kwfd3AfvB7U5e11D6W4j
9WT8JlvhRvsciEI3B5qQ/Vk0jDcjOxQsftBUFBzcA7gHhWlZwg0QkN6KImjxafVAmaSK4lcISMI2
64x1WEGwsAJDHJnlv6MnzDE2IvQadT3vrfOvUVa5MQkCOD2GGPSCj6M/BZEQPNNeesydCQNRhTOW
RY52tDhXob5PS6XEbrnOiag7IIUMMAz2iL3BfxA3vnqMWVSODGhQCz/T04tdkN+frvvb2UmeOcLU
71Wp28uznXeurrFOLfZ/GqvcC474NLs7nSSM/Jdou+Oqo03V50H+JBklLzbKWD3v7EAYxGPPOsnI
1L7ry69Wf4R4z8KbSsPVYcdaMmnNaw6ownwj5tsOUlPI0kucUTxol8L6jkaH8Wsp8U+h7/Dqouic
LX/zBc/zlxbpEH2iU97W6VZxI456Eu74oJaiBQ8iS7tAP1ExBLWuzSeGaiIifpXqnghcqzxw0s8r
gAbKaO4ZGBAzc5/ttDejjfrL22572NbsbO/GK9d0bKXNFWsz1tQvZI+B8MMI4nI4cvi+7Xh3rxM3
x//Ojr18rwTS6tVD1FF6mf5JIJHiSL7BgrwCXRnF+oI5fkkaQLRlalG5dCBWHIg+gbYPmg5QBbsr
4X7HnnNYY8BPMFl+UI9Z3bfx9+sPh4kn0OqaJGjb9geoe1JHBI+byw9ZE1A5NP222931k4fNpR0g
47of1L83w5sNTQkTqi8AlEVo2hMak855RUeOmxl8Nnt+qugz+nCOffl2xGTBNDlm0hO2cnDqVDMF
uUezfAi6Yq5Tao9XFytozADIjax1VA0BdEuMY+vuODtZZCpRi0GxqDL7pPbHNM5f+0hqlqzAhZL6
+GF7qd0ulOeG2u3mgu2ieG7MOvpkU69JYKxWKX/ExGMZQUxxb0XPZCsv6RJwP+qtvQNf0nlrpvas
ofNEkJdS470FSfy1Zdz+DbNaEUHoeVv04gW3V+bSoEoilYF0uM9tXFSZoio2DRquI4qKApUVEHPw
djF2tpowtsdssASCVo4oUQ/SliTiBDDQL2AL40XXvob1VhB37P3b32wsA1nc323GNQhsy5Wgm08i
x0yM9Qgh8tR+uznmchYUHRLa2WQUiSobtgMDLdkYY74NYSStnSoT4UI+ksYgye1zuhk3VZ8j/hDl
CgwyfNb+V9yL5m+yIjbMg2Qs8kucDxDSQTvTUztyBwuyk0ehsFpG05Oiz2mBmYFYQph3TiDfpg2r
XMqAv9inNwWI9Da1mIlKxdfYl6pEa3DAE10hnPaDPLZt2V6ZhjhDaAt8p5cqrPMagIzrmrGOUUdD
jJrvPHyQeqvoKcoezsnhJdsiZp4C3VZ+feTEpBIRlzudqzW1RSUauY/YuAykcTD85irIpMnDJpWE
bkh575MA5nO9Q0XxhxcJ/5NgCbDQAU4ZIJmXOk1D+JdDrLNUG+7P1h2ZkTuLGN4FAAjh49tzhqdm
zl4KrmgGc+WPsMbv1ijzeZxnhEs9sA0alyyeFvrjIdg448nCL/1P3RCOlj3Onvw1mQ5+9nZP/kQN
V3Dgoi5bQULG1/6dXc63NILQaFMHrNo22oIHsZ4yWutbLIJBa0sR/bIPnwf1dC73r/WCGOcfPhUX
W3+Q2hFNmZiVs0cwCDhbb/UjRZ5zy+6K0m8Yln5xF3AbEr9OwfdR7ousSbRpAkuEQ6aro9CbxY26
6TP8SUd4kTVjnV0NWUmOTEVBfR0PhObzuK6FpmLjlwRo20RVaZ79AR/jdbhbS4kSlVOuShHTLGDf
D6/lbM9tfVn03dWY6qYrPSXifdT1+8xZVOl2w+bnttoOE146mZAKC5NS4lFpXyxBCKuDm0r1l2Em
p10ZrtFIEGNav6So+M5XMp//kCf6/fEJDVmzBT03jg5/kxGeKdlIzbaQqsNkRr7kJo2KyCiXrurV
msn8L/CN/SFjS66LcMnRz2MgXw6jz8elTimsW4cVOgiEpfzrRRhOQNXTv0cnm9b2YG3j1eN2bRi/
TVV27J06FNqPtzyTd50K/14Tr3mF32Uo7VrhJmg5ZLBE7owRr9gqHXPYm1ycm9fkQBQ4Iq9rWkDd
Kz0//6ruaQNqxvg3eX/FghGiHkH7gNyuDm7w906TSf1F4lUhGNDo+qSdmkb+AMtPKdABGtWumWZX
jgdUuPVvIWKnwx0yE+5V9KFDu3UPUv3wgxNOTQodfiK/pXaFUeYTq6LaS1RSIlFT0eM7W2NY+N99
bzw9jJOy5HVV9w8l19Vy2mMX2sISUU6MvchhijxE2W32OXze/Az4A6cg/9L7mCj0LhfMqa9UI4Sl
YLVyzsYzUl6H8bePbqtplA60ztJZAsaqtNrfKl0KUO8xML1DXT2X4ZoPfrtO2+3aVtH5pLhTkHt3
sgMLG1w7xDSHLieIQ9mLIkQId/wiT6nS5Q9E3nUbStEaiwPar03fFlZTqo0o6n2JCl6LVIJUJ7eK
6/vt6kTwhcoVa7N8c1hJZAJPG/ajOY4qgn3ATm37xsdQ3h9lieIUb6g5z1dVHJbl6w0D3WPuoy0Z
A6Enjq+TpxW4kovaq15aSSFW2W6JFJqLpUAHaD8Gy8JNv9fx9dvJZrSMvv8InxXhAW/uYa8g9M/v
FkBBQ5aR69x45XYvIGNpNlmIDERWmbvehO/tHKzNnTQu6H8WEZl3NlSCC7rJ/lAEBMVfnKRZo+OM
iU4WPj0/t04znDGYjn6XCYQg6iZhgEzAT4HGtEa29JIqn/McmBpxZJHtWDCzfvZC+5NQOQAYNWEi
J9PIRygunJVTyuvfeLQwldkVkF5kCQt3DmFFO5XaLMUjagdBFS8JdQAgn3Z8WN2UABHOmhW1f0e5
SJqZriLAOwhnwgpLL++neRXLQbo0zXgMo3Up8/DtPr0xGBGTARsp4/A2a3657Wzcdh2NEWAhifRf
HfztdmApmrvMCPUiECL5ro+49P2bDj/0CMhh9RCxTMLEAR9qoEWDot2WASMS98NvjBG7oMHnjXuO
DIwLfN085d0Bdy/YwuYw7P/a7r0K0bdovnQPdsZdvxvOiVqwvGAystuv7VzA4uZ8FzVouc+1HXOD
bJxd12og0DhoAg8iyVVlxCYoUOMqESvcLV+c7ZwGXhOykKvKGKyVzL4V/RNCSlCXKzMS2NpYREFb
tty20ABE/VgLJbm8Pe0c6rA5C7rf+deeRStzCc9wgRxCrgoVcqukM+4qrlyDXr4L5UO74Y32aDHH
9mRwXnkq5dNw+b32VX2ZJ6Ojm38DEKzsNPy4GRWD0Upaf1muGE0B3ggqjZvbIHELVYMgxfrgT0T2
3GkZZlEFSD9nrhB7mgY2X+d7C+aEImNfcp00ZGU0haaxWiAsCOTY16+vmneHlVxCYOMXUYHdJLgK
mXkIFNZ3L1xEOJYYpXldRhYJ1cHUZRn9mnQ8kQhnpXsFhiNn0ISYRCY+YPnkjlIgxuo4lnPvnamu
y2pEbVeryjrsk6Vg4pGOWBQDXbZt8jBjMo8gI8TA/dyDVM23mRUr2qlpuXXaRXEdes0DtnwOxpQ9
MoGC25s8Q9ZmIR9qzQN3n0UPbna/4uO1Up+PWY+23KJ9kjOrfPGRMs2Ph4oji7UzNLQG53VzZSfQ
NY1mT2095xka2ZoNrpJCaidvkMSUcczdRgXwWbI+jlAW/vSavfo99SNf78AIMe9AO1S1uLsRmqxQ
2HYP3lNWIQtVMl1BcC2v2X7kNuu+TaI5+Hm1QgjNHAY7ZzuZt9XJnHCTGZtwFLvcrwiLdNd38CBn
8IKIwhWdu5cpuKTM+UtZQ7g+CjojV+pY1BgYF8Nhf1/SK2XkqpowUk2RVpP6NxrHDHCPb1VZ/Yn8
MzMQq4tmgq7jAxaYGpzZJVw3fqqAV/wOj8p+XeI3N/5Lks5MAYOvfvXrol0oqE4/dOmkfJH0rTEZ
h79S905QxlXVD+y3YAeiZ/anwUUBMsooM8I9D7aDrlGfnJDYLpGf+L8UWj3/fLAZ+UqsPQMM4sCu
ZkX2F9WMQtQn9lgJRV1di+kLTt3wJ6jsNzpORuFnfCf+e2RTXNEoPbDBpIqbmxNkO40/ZuEkJcUV
O9TutHeC8X7nnST6PlvANMAiVv1vx21CzTj3BlYCtO5WpJWPxEZqhNFZq2Y1t/ZEN7fOvpTPxz+j
Wf2EUfgIOojW9mBuna6C9hIC/H+PMPQA53DxcnXwrwYIFEyBiHJNNEatU2hqqmaaY6x4MC0RVXDo
AcqojX1Z3FLrQORyliaWRi8HY98JGiXKA8/vo39m8KQPkMiKmPdf3rXItT10ERevfMmLJT+SoO4F
OPZ8KonlJGhMQUYkzBc5HU7x6cLS2dxjRR24jVJvPXzm4kjZC+Up5qH/eJOvYIYOLq1/0bDuALUa
3ldVPInorrJZESlCIwlZ3QuuBFb7/ZQtCLyfiuYf5Cse5JbMhA/iTYXo0laLzgVW2xWhxP5FqU89
4iF2HEPdJUGUNJxv33LYGz5L9uDJVVlcfSWsD5S72OplJBj1bGgep6IdmlSnxFeDcT1s+ECOSBHX
NebwSH9RBuK6ixuosfx0blM6DNA1kZgANyLSF544MReLUYOeYXoPoTH5WgcuVVNDsM/Cb273Rvae
E7WR9ZuLMUktY/ROoWXpTx2QQEwHwxuRyL+e18rJZRfkk1XL8b45f4FL94C90P9imqcQmGDoTIyA
p90MOS/6z8+dJdlMJi1w1HStmqF5lo8bTOPIGuw+0yMVBT7LaLgbGhJPn7zYEdqipyfDfJmbbIDc
Wkhq9yFijLfbENBq8Iz3ymdyLSD+vCALcE6oxUTq7bDXfAQOVOVBDK0Qr37K+EuY256ymHmJRbKT
xHCsz9cpj+sJC9mhmJ3hXSQhv6Y8WwXhPp3IgyBl6VoHnjAYtnQaF4ucyriQdu62vxNj9A7ZPDh0
ffkwiRkY4gfgNZTT+sDNyyMkSbLXj72dtgH4VTdUr987h4rnvrmNrUlxDDE4/Z0+Mf3+0/MuTrPO
g1Z9o3wENi3f7+SWrdvGgHmYEC7BipiBpyQnc4dD/SpZzrBYNUd68MbYkTmQdzu9Xs5mj7+hfmEc
XUqa/54ExNYK6hzlRl1Ma29GllvorHhNdEgrcPIKKwEElHSCasMvLyRUh13sAA8ELUfYPb1CHvJy
pGoCzM15D/qXwKKg1K4Qta7x1+OUIqvK1hEvVvoTCw6TUGB2DWVdgnaue2CMby2z7I9NodOfV+Pz
wx8+QqE6tRjWLV6PQGO9E+gCX7ZQRpBAsCAQde/KrXP/qUPGLIgtyUVAorC6KyHsrOogJ+6yfckC
22Nm9f34LZr7ZNUMvtFLhMXzM2JuOayGwtkJhe85GFF2zhU5XAxBmP5IdB+k+vV5ot4PJHqdQvHy
VnTxlHTVoFTTjF4RziYtb8tDrkz1WiI085g1cCSywnUW49Oszh8fLfC9JOEpCTWbZX7/Y6pzr4RL
gHVTYD5kjtRhWCugD88VzxjfUfvljd2NCGloAVPgDkj7zvnWcjBL/453ADnXf72y6z1mrkQ0f3lA
jhAYjUjGgo5PJ9aQpRZvbwE4ifAnH6VrSt70QGBhRJSdmArij3W5Ru8HSYgiodf3wNj/iKC8f6bt
Dm4/7dKfYDEaxBxNlgv37wG6cqBP9nvUW01ys4qvSRSlPhenhmoqKQIydg60huP2Copamm1eqJXK
ISARlZW7B1Oyb9KDvMZn48nHKOxet3xJxC+Ijbek2jHxCQQgMiu1U4rKNfN9aHh/Mtxbts+pds0b
lgf0SqtvNIYJ6F6gvIIWWBfLcrZxO9kjkEWdzFj2rJqo5Cgwts2yTwpQUG/0Ohib0B/kWb+D3kB8
wxme3QeOabbBjH8lIF8NYeQGLs+R6HxoE9j2KawTt33DThzjjpUDTW7kaN/USrONn3FHFJpCL7dc
DFvFFqXka+uUDfwAimM6ZA2gDWXwi5Nsdu4m7Ob4WSYhtogdjinR8CrXmfSvE/wOvX+8Ml/mnyxs
qZpolNvFxLRYH/3BVk1akuAPSuocPRXoBNQnlas6U5o7DfpSDPy3m3iJao2qUDMLb4fJLamtk//e
ck71IF9kfH5ccfilktmRMHBaosyzyj3C3H5+jKPSZvGDGoi8MF3dJ90OOcptUAWaE8MlwGlBbGjx
hsGQOiqoWot9WC5lyunet7up7ITzEsJ+YpCJ/ylVfMefHlF+uSpzS8ADPFpeGQ35yk1Na8iu3nwU
X/TTXvLMaYf6OUgC9znxk/xTF8VGRII2ihVC3Lp9X/JgtRT1PkL6eMpq7OBvGyhiJeUHbgAWusdq
sdApZRIY2V0qiDpVE911oaQdhWAU5+mP18wDMpJT5GpE+JEJHiTXmgc4LqnhfaBSzjG0De7KB+Wh
/VsyXO9SYBvl+kyZVy7pwKSJ8NoMZsryvG50w6O9g14YVcYKZSA0GNU3n5/shs87tfCsdeRlHol1
hF/aKbIOQcsyKBR4EZBRRGMvN/JE5xjCSzHCutgWJiz9rk54sOM0jN7Vi3mPHSF6BAg25jy4GnhQ
Vp5GZk+1OyrP2mdZ05d5g9h5+LtXOt1qbha3tGqQid8TLk4FBth3nU5nJu4VzcLBiPSgH0vF5aME
PQpFU2vgGsOaXsboo3gs9MlpN792ddChkS3o1yv9ji10tvHAdCHmFJm6OfKA59WNxM1WwQ8WLuKv
EU8Ah7i7u6kil761NKTX28wtYWuydDlOKbY6xofEiFHLCJ3g79CskO0MzemeDP+2OR2ycpTAe0vs
1ukAruTRmdRbxDXe7Thcp//hGm2rI+7TjKwOBxuxZGptkA5hVyogk6KSM8hEMzWiwslA3owPKQZL
YcrkfkAZXra5y4LAa6OfpElbYJjfR/MVLhhSFtGGv764RYJyeIllpNYBWGGxSkK5LKk2AQJ8j+c1
b4GQ/DiHrejziur8xCBZ4LJFlGMcW2Ky2ohDYaVCvtY2UvJsv+PQNbRLTZcZsRfRkfjQgpuQKOWo
bkRbnu9aKHQVjbQWUktQ8VYN38jcKLrswjL3yGEP2ldhintvvfNnQ/0mJlycRXT+o9/PsLTOTwDS
FPVb/Dsl7bk25VvUqQtjrMvUQaNztsWrSy6W3UoqcNR/0SO6TmaO3sNTd3bxctx7BnmVREtLa5Et
cc1cyPZSMGLb7M1RsWTw29YXdBY2NJ1Ff0KGoTPY9nrQRaPQyuaha4XWkrYdNzbh4uCZ2jajTazX
Z8Gj+hUdS8zxc8udHXnN/0k4AEyLkq4Y4/z3G4moGOznNrL8Rnt4YnNStifB4xuffulRFB1bU9zf
4ShtV5yBGgjPuLaGFhehJe8kEPDDLh9QH+DxloZbNcsbsi2j8cRaTdHTCD4BvJU52ndQPHUmKuZk
XPvfVowlS5eTJ+t02NoB+2D/biDXHBLw/4lXU8OntztY1WMB3Dqwp40ekF615JeyJGcDkrqNzjqt
JGKitlEAOn+OP+FGOr5p06YK7i8WvwZ7LYKQbL5lruG5xAT+kA+y7ViicDTrLAJZALaJ1tVElwRC
JIAL5GeCzQHfVqehl4twtLue5u4yf4JCBiW3EO8WIMwfrLVvTepKboh7RKl/2E3CoUODvknTNNnK
h0xqf7XU3OpgI7nTELVldvC36JVC0KoYkte0J6eUWk7Hpf12W2cc11Chs2zTodXlZlD198chF3C6
bWbZunX5f2a0gt/a7l/WY8mMNgh7LHgpg7r+OuAXIoLtANRoiZRLynNcyMGTEiMGccOMIF4ULZOo
3d5TUcQ3Ral+/Zx+3Uv28SuOyJYD7VV/UBAsUCFSz1CKsjtuyxAPZhfOOy8INNd/IM/2MaqZlBnm
ymQr1TBI8tv/YHLadTqM8QVEMm+mjkm6BGMn4KYHerrAxR6F0c7NP1tHWOEexBTt4vtmA5U/ly6x
i4G7/P4fMMqZ1psewJXq4pyf4E/GpgctJkj/lK8yAfKVBXaaBNOKl7BOsN3cYXvRtCRZ/SaM3Jnl
/9OVR+E3bil0SQlNS3AFKdkEfILAppqtWM1nvh5uXFq5loZCT7UpkZzFIGhEeAkAJnC0sq10ON5S
PDE2MyPvw/mvhwlS48k9D+CJl/E9qAnV+4qzpCQxkrvDAj7eMR7ot0nsmM6psCzMOkXpJGd8RY9u
dhKdwWMtJnaUNssTvaauXVzO39fOt00macQd4Dk1A4TeqbQSnfC10awzjk1E64OygZbAaQMudVqW
FSZP6JfWp+c90tWldfg4KMDPZUvBYWEcDxRfNzD5U2vWJSdc+vYTB2CTORtH5ggI4V+IGjj2nnHl
AS35Of/N9jkXlZuvo8B73oezZSJRUl7b48b2I3OfEoBSrJjTH4T0iXb7cq5JiO1YP+1IAe4UeU3U
czzpVJhUCoQ4jco9JnXP25bknqQgIxBmbXETFB4Q9E0b/ctGHtXH3HQ88JSSoAb6e1zUI6nUqbm0
Cu/y/HWT74vsWnBy8T0p//P1W0Z0jUPz2vdL30xJ2gTv7pOJIj8Ju/kbe5HI527x3L09el8tOMpt
SIETBZtzPP5jAJzJwZ99ktfCCJJSqc5hRzR2X0hX/jNK8AMWVbGrQr0AO1AxX2yupxYmd3AzQ+vU
wj0juuKlbccOWhxTxOtVdCELNGVW4JWCznxPM+eW5Rgnq6nq7kQagnQVCveGuKxxf50PKMGXMLu0
ud/o7MiEMQlLaSe3ATUFDrIBi+yHAzaM9LFhTnqm1Brughg6/wnqEXr/eUC8qgQ60l0yBoeRNS9u
qKCNYCFwNQPCAnn1yMVS6ws6puU4MRTd3RANYaVr6kBuOvS5tqsgDT5t07iAqzgCHwBxmy/8T1se
Vf1zy7RLfeDze4NiSKM6+yVn4DWSUAo32ICl3uv+PARapbyRvBsooN9jTwRDRmY9VDnl231WXojk
jAGre71jYR3M3Ag0HA/cIjpSdy8isSyQgTlK9M0Zpb3mAOJ87e5wIDOvNA90YrD+PeDJqfHc2+5F
EUFsaRTVWqXBUA9yM/v8QBC2xSHOL2qgnWh4wYKNLT90kzeEE7VdK1UTJOoh1GOGWUasE8CXnSzH
7gRJ0MN5ojjGfJ3zpZ/k2duk16xNAbgg0rEM0bctJHHwNjEba/Rd293dofsFVFv/4WP2jklxwhPy
aknA4w8TP43MwT9NfBmvdjrpTceBG4hUb8rW1uxEsOG0l0J5+i1pFS7uFADFedmRAFvKvQ8o3png
hyQr3EOiORd90sfifwhkJj62owvFpHe6RUncYqSSa2GCudSZBCffD09dvj17W2gVg5bWoyXUyzf7
+9XElSuWt/ZiwGplxX/T11w9m5/qIg9sGqU6JhyOb7gK8gC16wmZQQl1nid2Q4NMtiF989vZ9oA0
H19AsFHg6o1o60h9EmYDvI/SnjJFsXplitdUIaoUMKYltYScOQCla6L4I9kvHZ+mKdAQUIPCoq7+
Asp1X1SlFsV80EEDN1aEbRO8Ms5bklCKyuHXsB/G2M9BQSDGH5dWdJrJVc4QTKsvbH5rJ72Ov4jG
1a0N6uIOxNgbrO8LJavkkGz/2goMRz+FbSfec20cRV62g+GtpBuZ6M3wU2FOJI4fi/RcR9UjkQwb
LB71yGJ1WsSTMADz85HssjTgEKukcT0IJuljkemdIId+063iCpfSJyMuq3vI6TTFRekLRYKNpMPO
4KaY8Z9YfJE+VfI3c1HE9efLx7jFjKWTIB8fBn/WKsrFkw3cqYQX57ajGBm0HKxiZ5Jii1Zksc0p
jiS4xCYgILaCN/U4r8SueQJzJqvvd/ziRhVzrYZfwqjyGAIfB0J5A+yTl4N/7HGHEzP8ErEVJdU7
T0A4pXH1aSWlhIcHoobPpVrbBWbbNZZ+itPu9aU1DnUjEUjFyyQZ+D/wyQi18Pqy0BEVv7rTfyUp
oSDsYFV3MMSjQCW8wqODLznyiK7s3pmCfP7ihkUXw/vLOj6EBhGXfYIt0MXP0VU1DKgRcbxRGb3b
4owW/nx5HdRBxQEnSmQzvvqUd13kbhoeLwNRWiU2T4N+yaY8IASqJbqvENwQEnVW/p6ZcUJ6mf/n
8QSQQ3QYxMrgmtOpQeEz5MbMOPr123uyajkzPHfuiZUUIqlQjU1ogf5k5bWsG6ar67qoxLvtH/9X
4gF2VAnwGUGcPuS8MpKzF70Dh7HS+OnRFaBkQYQ5ct0R2OLLrRM4XaI3gcZ0wDdBcseAzXPr4yfM
y2HAolMusezTLdQOLZAS07TcLP94KLKvxGKSMDLJQfdRN381jrGT+DIm6YFb03nu//P63tbjy+iJ
EMa+dw1v4WazUJxYpHOLyuTWVK89Ofpvrd4bM1DD39LZWGjKZrcHfU0DqQZx/r3c4Tx8YVYPbsRP
Ir2/VA+zGyztFE9pi9YYRM+4GR0wKT9Nul/9NKTun68N4YJp0EzjaKIGTDaykEAsF3+NwCxqauRj
Umv+mdd1V6hOxBCWAFJWB/DwZRpZWRqq3hLbdfZY3S7uftEauyN2G+Tmu4xk/BB2LmI82ocQRvUP
ReZHFvYjEQhLKsTe2xg4uXfKLlQx3+5upzG6iYRBKYy2BZPCY0d+hKOzLWc7jH4ugU0hMMxWnt7X
ZQH8K5hfhMHkDQJZyxz5sp36rXEI0LPgPoM6HLP7NkPRCGpdIbwp67H5KXd7/TFtrqJF4YIJPYJj
E6sp3KFDjACmt8eoAbMc4ObS2bdZ/+bqYxoSQR28ZPwKkMFOEmZ2EHHs9ydTbAuwlQR4AGX4l4+7
SGInxUFvmJeJgaWBUlReaGwxRwuAM8RBJRYs2XOuLC1b67cOM6ZjEbhyamYWwbdaP5+3tI2M8I6a
ilfxjDiTR284rBmlIN57804wkqfqhkNZub1wzZEH1WWpg1xywGvDO+amyHWvA1gjDTCgaucSLmVc
Omm5NYMapYHs92Md9AakkQYQNG8jMDKYYk15ltHAipum7ghqRtrZCyjnFAm0Feq+3CdtGR5QW18S
AawdNluZsRpTT/SSIz6XW1wxII0V+58y1EprppD4L31EUpkNJUdTk2phKzwTHcMd7MszWLltnLZE
ppVXtzRqdTSb6F+1pAm1wVRi7I5wz+m1T2u0tEBYHqXaYE5LLE+yd44/WJ3UT8YdZPKN0hB6MOLx
7vUdHOnLA5FxwB6tyBNdJGQksflB4zL9vZwRHTsq0HO3vu9iwfIOyfO/ygMqoYoieQQ4lBt9GMdd
q3cfonENEONK5XLiLlZKNYseLv3kVlkCXDeG9zRRTwQ/t0IF/UwclSjC2cwdnBmxpEcC1QvvV9NE
Oyy0hIjLBDoB7AlHsYZhnC3R3PtO95hUsDTtI4YjcGJ/FdY5D717IgHSaBQdFd/pW08lrszE4S5h
PQY79z2jI0LR6N0sJMtwBgI/jfgrhQLy+EKQDeSSiSazwU3Jw+PiKNf3obb9jR85tkK7zcjLSmDx
kOZvzcLnxH7scC4JIf0jdiMPOa98c03BmKE87fQESRDMQfPsre1pzZGRdyGwGwNQupUpdprrpbQg
ZmlEaqLx3qzin4IrOWXAvoXLqT0mR+S1BKkY8RSt5hW0OjSrFzL4jp+EhyY3kkSIeUwWMRrrwxQH
RXQPJQNzD8aA/plg0lL+397ez/F0c8mqHMezbwRx4KmiCr7O0KAltmiAKMllNwmtufbXJU6r8SPI
BW8zzPffPKnNOmtgPh5Z2r1+MYtI0GTjSRLs7xKdvyOr/xdGgv7Q7+GsNHm6yiL2CYDVaYNfcO49
Bi21ZbIZUR2hgGweA1Nu4eXez+APUCu6X4SknxlBeXb/0PF8wjz8Im5VNZ0T/4UsFvsTq1wH7uTH
jUQwPPhidvHyUaLIStBIe4Rxcf/8lV3KxC06SFY3q0mlWpiOnkzIjlEVUOPYfIKE4ZLB/xfIVKKM
gMIN4EYwHKsdMwfwWZ6gYz1Mne8GDE45MexpzUovSNGmItJ94M9eZEnNXPRmTmve8dZZgwRJ5mMu
d++2SULQKOA2P0bXCzjrOO7EluP3bsHwQawcls6ihtbewH4rhlTQVRBr3wUTqxr86Z3ym4IhxKjO
dtxoBfu11+wN2xm2rojNh0NrY2RIvoyCx9MlyEM+usst1LFZ1AEOmsiOKh8uALi0HyUcbb0twcEk
85zVRfQHmkVfufI6a2eZNNYl8MMOBt2hEmGWlzqPPn6xH6i8zZpwZp3x4IBny9dd+GLqRZAqqcdl
qFkFQDzhh24C6Gg3b8LnoH5MHPK9eQ4cTDc9zITUOf4bkH0OJzTaTQiGJdS1xd2EPRRM5TVUgDzZ
IOll0KkgdROGX3vjAXBAJBMcGYYp8/37N7j94FfinqyQv2fwVEBw1Ha14v6nuJQZ1U1/9I/BBVoH
6yaRtul1/5k/qhTgbtdbKSb68wI5jxNFlO0+zSnyMEziGj+ucgwMPWeYWJeFzfwzQRkq2WJVS/8B
a4CLUgGtPoWm2aFkm/yUh1dpPXU5MY+dMDtCLKmGioj4X2oEn2s8yPS3nzUBb1poZzZq2MrWKG+v
NS1zZgsOog7n2b6IjaKhcokRmNbUkE3Zp4+NEc1mWXmuj6h/lC3rZqgNRh2r4yIgJpyIynC4Eo1y
zjyhvKB0ujgI+LbL9lx7adWxHaqr4P4rszjPMM7qHNY63sbAsUKmrYOcT7rvbaRLKHR38dnjl5LG
j723AcB3S2Y6sWsuHLvRkuh4jnLuo0575CWwXT1TLO/lOuuHzIqEuQOqo8vciTARET2V7lDC6dN5
D6dm8fHou7bE757Er7HcKkonjY+k5kCEyNTvMK3s/aVTlU5HQnBL6P54MyxkFhcHwOB5kIfwMUsr
hp6SLNpKIM4bHVNOiSy3A0UD8u4BSuy1gx14I1R0CsDPP1tUVEidCK+CczJ/sJ83duMEk0CuYopg
OMN60fN3BrxRjwswq5fNZmjHUquOSLElZwXekpAMvp756NvB/Te1RqzZV2fYI4xts+Njsfpq9chp
BLm0BmMK17sOOjg9kiYo9VT7Wnbffj7eBtmi8NPoIeCm/l7vXX0aOtQ5AboXxBA+PHJPv/DeEwbs
ttxZcBb/bKgVYgr0E347yz4rbwk0/YvBVOPR4ogxFd01Whco2zRKH8hwdx52OmCm1zuDujx5+Gl9
A8XNoJFQiWn2fqZ4X/JLQpDuX4mkJpbj1Yge8PP4hTiADbBSMkjbYCT+DPp0Ri6lUMl4Qng/nVr6
vXM88QLGbnO6fzOmpR5K9xS3yow8zN72BOAmrN27DB/CsMZ05NDicot6CzEaHX+vejcY52uW3SiO
jElwNZbDJwYukCeR6GMzHLM2SvkuG+Nr2kjwRqeQJFMRHKnBSjQP3vxJZgu3UGH6WZ6Ib9KNvdge
LPKljrJOdCZDazQtZW62KsEIvY3Un3PDNwFaQ09TZ5MNxxCO7n44ZOlX19293wuMZlOAEISf0ql4
PstkcKMAd9Scpkxb5DF4a6RCh/Mj9YiuCDa2jKhRQF10xZlagDfZ/5KUNBHlqVSY0qyCSzAYqftf
yY0HXxqu4fYhGRRr0/xN4M6DKZffo+R1MGHTdhfrTQn6kXT+lYyLuSfT8z+kLaXQfUrZOZCv/6rm
hdfy96kU9xUntguFWEfaO02nArHFDApu3ylUZ3V5WFFh4V+jbYcnj6N4VyZ1uHc1AQTXYV+IaDAO
+jOYxu4vWB80x403EyyVthOto5nxfUwQ5NK1YJrRtfq2m+r1eKwadjkmujCZ7iwyYFNC+iucY7Rv
IVoWF8fNA9SvXYtuG4i1pyfnhZeXM0COQ85LR2rnHUUyBBJC2dMsWkJjFkQGOdIJVaPXnrPr88Af
DjwaGm22o9AoGndIF/mvrgQjWQez5C2QPs1lxOJSWCvdMAhUIdjtbwAzmOMfM7jtvfN2a2zIjS0U
MRrw5mf7UNAHPE0uQ4K0NVolNqz45oPjT0LUT69VgdND/JWuH7BQhch45H66KafcmbRrNwtB/euX
eBGw9nuoK7K61Bhw+gcPGlNbaWV+Lit7WzYkc+n/8LwHv5cJpccveaDOUPdB4KYiZBJKTaXTBobH
FzK+gCCX0QjcPtMYXE/+KhXnnyhlybh7IqGAL+1qmFTb0NV7gFAFmgwPqKcaRY4rTy+eTwP0L8nl
CTVnQGKsY8kuRa2tKHTwgw8e3o38VhkoFxxTTGPTi+j7oKQy4ODOS3V+x6a6dP8j2WV8IoUy4II+
hZ7EfWcEhqpVTKeLja/RwKkz8ZJGw/8D+qvnpcKXFuRQyaUPklIJQ5Wh4mioWAY8MNWRqZI8D+iS
/Kd/+/NMlPtHou/16g7WFFcJl7daPpsX9QOxckZ0PbZRDL8y3k6bgNdaYBNm32qP16c9EiKF4EDQ
/G+ApOZhbFpr0QSqWAqv29aBnQ7DqC3A8kTjCtM4hQKffk8xjI1OQGoUtVwjd7y/ODnL9ZO4xTMW
AYIefD1OctCDbaA45K/L/eHNAQjP0FzQlbpU/kwHDcbKzBM3psr0SELDl1krBm29DqU2oAte47v8
Pk5fRUtTjq+VKxSlWfguPriCpJzT2h+b9ZSEs2FrCn5cvCgON9nq8/tOv3X+TbvADQZD6FFpeeRp
QCEdxKKRef/7xjGVIwkaesBflAwYSQizcuXYk8QmRcrWKwRZ/TtN/HvBU5S76amiVrTkVQkYlKoG
KWInUbKKSYI9TWgDl7xFOMBLF6OuqxgVmCvooI583AdnmXMjEE2san3LJ+8SvjJQM1U80RC6Du3j
d8mud7ipeBpDOdOoZkBqIpV2xHOHgjlkQyfMSCqbKHyg0sY3a3y8yE+4FsIYTiM7jlWimrhr20YV
V4QsGDu6e5jJzyXQx6R3VqaeHnbkv955P1OefoI8MGwO7Vc3OMOQBOm/vgx+A41mmk+kAwCW75fd
aF/3nTNx3re67Y/XjoRFk7f2LZutEdjHcPkyRNwEOTYAe8kpvSkTPXJzBM4g6W8VKZddn8NQF8a4
boksqehzLFHp0e8/JCJqwWAA+1B5rHpu57gf2Hvu5dEVXurSpu/8C8zzGmdJlVDRk9Yzpo5m09HK
+8yBkUAji5onJggINuAxmavuPE5z85IoNZufdZUET9FuYQVhaF4m1k7c+ACWCI7fAjjlq/eHeS2q
cfCvxpq0IitPK4QuYyUBILOQh+rQAlqhQR1gHSWnGtnitq26aX7KC3GIxD7TByj8pIBnNGEBBc+6
dT6QOumB1SRoMG7vMzp4k3gb/4/o8XXALUiYY2fDmD2Xi4F4mKR6voV0dfZab78lTs7+GEViCa3O
VjsnotKueHGzR3zMA9uBt9uaPCqULqHvmNhAbhuB5mzmUEMQqrB9TxCCBaXTpy9vWBBoDdhCKRtG
eWNO3zelPTle0Vaq5GE3C5DE4yDzTxrjYv/Bl0nz3LNCPnSjATCocikKV6pamAqOm1IiVk5jen6o
iTOj7ZzUjZRVjGBzaL9clR3UOooz6ZhJc80kRhNmqueFk00svJa0nd/11kbsjO+nTJXx7+6Pvv5h
Sa1AdBT4Esv0N/VNFULxvT0azUomgIvqY5wIKX8TZRHDT9ouNs3d2oGz7NKy52ISfbS3FmVrbrtl
CGLDLxy+HhTYJyboU2DjWAxVcllh7071ZTeVrWIGCDBgX8e0seDFPILh9LeBIAM0RYjOQRLFwcmC
ErzkY62Xp9xcyEiKh5z7ie+oAihG6Wo4a2u05zJF1HT+ug1KVOrkvbmMMmB1Rt1C0ddjSQjWfyPx
q/WhoncZj5vsS+ZaaEYkNYkTJua9hVJadu07AXLIDqjA8W47TVgOzsd/Z07DvSsAFnkUTkBKRVWB
x3sgsUGni2pQxNqwcNsiGuLYIebjqt34NcIP5TUqlAyOAQa3o4XGIJsZYrB6w93DD4G927xo+FPe
yw5cdIIg8bMlkit7Q3bUeijl3H+HSU+say0rRyhc4hPsIluJA6ZGgGmAvnwHV2wFryDOhEj9kg20
l1Nl+MR90UqTCxoNI/KD5axk45BlpgDHjn1NOxddjPT7Ka8X+dOOIr1Gb+eMUZxdWtKF6pn+K/KQ
nuWq2c/fQ/CQKnH0CpfkHS/9OgrYPH5AKepHyICS61y0c382lT/R2NHiGxgFAcUn51uw1rjO9rxO
DzQq6QY4/CBeWIBMoPPEpqr1HXoKcH/Wxb+XMaFxeP9pbNP4447S4ga38z3B2/khD8jhGPcKxZSQ
Ohsvf1I7eHzQ2J1EqUbMRHUk22FrsaEFdgraYIYo7qfbaHjjhOXgBH40VE0jidrYAXJNljxcCOff
/5NNzProR04AVb+NYr4xVD27GrPcy3WRoh7BYqE43IsSkwCAqhKB1PweNq85WpT3EvjyW51g+Lwn
7XiHxR2H7BqjMpfGy+JNdN+5jtk5jRkk0hRmsGObUUF7+7Y9Fg1XBxbDRd/uFzniMwu6lVFWXC3S
y/ne1p/sJJJNWeqxIV5Os9nTYfviH8roJ4FEJ2VxYFJEE2c1i3bV1vvdrX8rYDixrfkYPKWhywoo
xCOiAEC7HZk1cK9GnwZp7QbVwFUSd511S72rdZpwg2TDA2eerPGjw2BNuG+vkHcG/OMcJu0kFLFq
rAaED5Go9m5WIhFMjXAIG1rwC/OfLhPtQ0MrNC1lYrq9a47D0nhOvQXDqMPiJYK8z3w10fZcE1Y2
UYbjC3/elom+WygoMLEGS3vj4jbB9CS0r3jpGjgO3cTWguvenpIF5Ll77UVaVZIEWgiA/ECJrPgD
4smGoxxcXmRE8NtSJgnkzfo2nKS/an8cPPnduw1hq4U3mUTxckEtZX4jHBVT4TxuvCBHGUGEklCM
nw2q43ccovrdRDiq8qwcG2RNrmJoyycbr4BO7iBE8a29JWZiktAhvIScAyftE3WYl348g+8yQh5j
XsYVq2L9gYU45mQJyiIbscPE8ic+j51MmKmgBmDfysNewqxeTRZoiYBvAulPzDGq8i91SVNEi6/H
VtzXYxP8R6CoOIvIOOOYdnxMBOTtt7zXIbRFCegTZl+HLM8As0E99DUs0U1tv2bGJRM8z5HZ3sJg
j+mj+yW9VzdxM9276hVZa0f9A4E+1FgTyRXd5LBpQRnQLUehB87hJUiZCtpR3tXwJ9jVPUHOhosO
UL6pt8G8QPeigkn1WGA7LRAUrgA/4NG28Yrs48JlGaenVCyWjq+B1xghP2+RHXZcGR3ANmQ7f1GU
9/g3YTbLLmEqlPFxFmoobNaCvFOmDWGKz6DkhxPx/+n/x0eJd//WIOLdZv9VXEtV3i87hPcaROpI
FOJEPIijzOT2zbsEXznOhuooABpLuYW0SBx8WKvpAmLg7+nahOo8ahIUK8CuxWtXn1Yl/V/FM7Ue
8MsZ6Fcw7LY3SzqPBet36Opsk0meRNmDuVxvcjmRGUU4A6XJHmMoFi1fWueLpzAzLqP+/MiYDK+s
BvQpPtPkgBkG+zGUNh1NOV4kinLZ4lT0+GuUJV/180pC9+NOdUeZQZf/BNrCA9L1QnQCM3X4emJ1
yGrTRHYpLYZ3Evgv2iHguXqJbTwFjBROmnKDhKxVusLEd6fNoHX6LcBPEATkPU1BlBSMJct66bi9
vvc8rUy4NNFAJyCpFsP4T+j2Alvk+7OMlph0hW3Ndot3dHr7q2pA4x7JtRSVmB6AmFyh3fCq3tct
nGGOi8pm+Wu4bDySm9bxUDHWgv+0ee1t0ShPJbJbvnCNNxnBhf2sgMcdPTgUDYOjILiiWLpfVf+M
7gBmTMiWpPL/xGklocVdueR6Yqaa38WhViP8EvsT4vdZuEBrE+NNrUL6TYKQVoW+7mdStRfWUFUG
zwOa+1eUCHv06BE7nu5BhFpx9s/BSP0ckjhSSijdj+fvpnKOQATjYi9uXJU4cZDPqc3vp/Wl955I
vhHlQ7m62EN9n3DLjMvalIFCcl4hfG8qV8tUQO6vQ3Wpv3x9u1mUtjpA2t0sDmdhAnp0N9rB8k4W
xzAOc/n7GqLKbkeYi/9uZ47a0OnFUZEbz8w2f+utx9k8hqAzfG17jX9mgjrMMGdhWF7ekT9kWsZg
Rm0xtHPnxXaiTEPWVdD4oq0VzVGsQ3cnN5xe8zolSWBHqHa/fuE7hBoCfnvMzBPgQehTeIwVd7U7
WicJrL55DyQhGZ0HSBGq/5RjWDVI/Zo7OmSG0Cjmxjr/jASa5gV9bG6VVEKJg0NiVbm7VVcYE99s
nrdwuAiPNWJgX/W5JedovZdG/5ddMWJVsHUY4KPkwgv5tGxsX7grfSJW0s0bpTFP0k6qlUm5BYhD
/2skGC1cT7jiCQcpW8MT+z6g4FBgE0sbHV3RKTMzgHmKBsSd6FfOHjyYfBOnTxVR3rDfGr9oUoXA
8G210aHmnQwiFonXd5pR+lZJY+gY76ddK48hz5ZuxAMz0oElBDaDA8VGod4eA/+1M3EnbrF7GXHn
y0HAj9AhQlsktI5CY3nBS9MB2uzz2gTLlGBjZbwI9aR2OWlWOpPrfuYANeUgiEtMJ3UvMeoxiwQh
/FQkZaNIKHc8rLzHF4EjrAeo8Ms+D+NI3Ldl5U9BHB04mxc69lPIhJ+PHAiCe1j0kp1piOT6ucry
JfylF384kRQtVXRuuOPDwKKvvAEmVDOJ8znpllxSBq4eYMA3fEZUYKhGVGmyvczhHHsjJX5wgy2x
sNgL10Y8oMqEUIFv7vnVkEkLeWiLmM/fGplQ82f2nuQZ2wt9pVVgQhss6QEdl2k2TvCrS+K+mqIA
iMdRvWsP/bkg1d8LeJXbLZjE8BCvDfMCcpiQzHHzj8S+svozIUAmAATFuGM1qXJxybBFp1EIkHXm
1terbGSAWw2DTyfJFVspxL9vGPuOFSU9hLXaVsWqDul7IgIZR9fsxeFdyes4XYxalvJSG+7YjOxz
diqMC7MBF3RJ5KNAAshp2c8jczhHlYMIJm26pH6o+i/Qs1DJ0XqjhKtMvkcMId+DzTKIYf47ZDgY
GcD3/NDPneR8rlHvBwfLSjCJQNqxlZ/d+DxU3w6fzoZXzFZ3QxhWAabva48dY0/1cIhnR2m0jO7e
dISe9kwwH4MqpoJLYzMlPSO0g230mdP5nkvyeKsXTZxdGW3o7xnkhbTX5ulQmTXjchArgpXdqMsP
FBpGNM4naOZbMoZOT6cyvhAI+PAOVGrsm76CpKA6sfo//4DG62ofcCIdjq9XZ1A1Qhd8G6CwUN0U
tIZV/wPOXSj0+d1ZbaOvWOXAmaOTW86QzPjROg9SUhu7I+D6TKslMYUTeoxB0/Mph3GmSnkJFxog
kNsSuo9qlGeXR7fuhaPu+HlDsJv406vVan3uVxXP0dJodmacMQ/VYSWaZuH5V6DeLZJSMCb+6lxL
yythgIZBNGSVhC+SaqTFoO8TZgE0yRpWzNp27975u0Pp//eTMfI6NT6om0ZGD5k2LXPcRp2T+VVD
DWjo2Yj73J2OPwqWBYisTMwwLD7INJO/wm8OngzPUz+nYVXY1As0oHUyxjFuNjZXNd/VHb4nPNiV
5qYuYHQCuYiwyRl8FcL1/oq4LHVEpo50sFjPVrfnFD0fyl01Z4w5XEA3ePTwB7FX2zggIOGc3DCG
BlAfoV7S24gyFTYNmFje/hLjZVMlREHgKlMRtnaR01hZw0yO6yRKTvAZuwNirG8VKclfSmwyIhNQ
cc9CDbUGhw02DtEYVTEBTa6yXS+pmR77z4nFX1+pP8vo6QyVAb4tSpdEqCGJDLaOA2CeOWFEGsoE
AtWlR44jAPz+f64rdtSF0LanRiqpMhu1bAP/KG0cmc0j5UQOUcmYWvkOou7Fvt/mRcLzkrX4vBbo
dVhFGsthCTMcBgYV98rJKO4n0DIF54wg02s/0JoCqxbn0pgouB0IpfpjM9chD6laLCglPzVGQ2/Q
bWihTGNU3YV9mulBc8RKtcYh1E9PrZCF2c0O+DMaxkt1wApLav8uqP8wvrOhcN+ZMI9LjvaCbKuz
5XBAG5ZJQcSaOp7uOgPMLLIjdXR9wWEx9xad9cyUe0Fc1iBXhcgbYmxhpv+TqjQ8Wbl0ZT6WUWE+
v6N8+cOuGFQFTFXB+Jj3SIVnsfWY7EDGKLOMc/5pNwVR8F/C8EcOcuXh+GcJQcswKqPaNCTCK/OZ
2uSi6NA0Rpm0x4sgGH5wsomlERIByCBBrCZx5Oo1Nm079b0SbO2AW1KW83B8mp4hFWae1SOyPKuq
DMCQHLJqYl/wJV4VHcbIu7JFIBJFPG0x1PbiM4AAbjI1VQ2pQ0jTlWGtKZTrCt/NRO3MLhjQiP0t
QLEc1S7ZWjchEm/GVAElLYAqDUJF1w2xen5bTLOV6Upur07mmiBNQxB+bIC+1i9udlv+031SmAh5
oV+9XYbDdHqAa4T7xVdhk/J6fuJ1xKAyLwWHyLNWeIpedNOfgfdph/0fCp4kV/FxKQmqLwJzx3si
T5gCEmrTYX9bBMHYPlYkwJS1VpU+p+/NQb6idvA6tTI/4BxwlyImkNyqZ/HSJkQ9Dm4TDSPWq//D
dLCgK5b96Es/jOgsms6GrWuJjwIFGFn6auu6EFps+M9XZWv9CMj6iHJMAf/1keWi8DG76rmYKoN4
kPA8NV3PnDL/rY4dy/km/e3hEBvm2W6cVu48CEJOfMnBaLPWDWtMwImgjzTv20Ouegq0KxqPmsN3
WixaGaq7LFieJbAG7CokjewBZOq9Fumz8QAeFGUEQDjL59g/+pYQWyVHLUCWx6vYidX5/b9YCqz3
30reDG03+lZXd2Q7CK7eotrdhadLUwxIhe1sOcjhY7IMxR5iFwQ/tAb9IQfAI0Vo3F4jjtbWvxFF
z1785zqtELpG1axvhKAj2JonMWaQdyiMC0ENYJVVlX6ZvioXeK86or4iSzDNL2WrDFeZXTR+xLX2
WwgwcDeOm6368pejxLGxVxYWEu8FJlEIiT2yIVttnSpQL4i5oPTzbHLagLzaRKo/aZXNOPomoARv
ejy1iPRuWwMkTlHh4W8Jj6jQ9Oi1uevjSVnT9cMezlnQTYYyNH4DAaRk2h9jjsB1YJ3tY+M1UfKn
rJ5wapF48avYYP4KBjWv8EUWgaoAlUAc1qqDKyeeJ7YaOm9LE7+4shdrfSsoVLMciqshG5aOAyTb
STSKHT2OHsS6y3xfOypYWLfl53rwQ57x0KygNHo6m26hX07LHLZZrQJ1ctb2D3wZWejZIll/Ta6F
JwCpYPpVQdms/FH7vVT2bPuwU+uxrlM1kFXYFN2w3oTgHlzrb7CdsOphJlWBKgHUO7pFymIeoIYe
NfSFf0r7dGPqbX5sSArNOMzUD+5pOOG/n0FaU7AbLvb1xDPiw8XSz7OsUXJ0BgvCO8P/a1EZeAbx
GosdKQbPQtDQAPg+b41Ute6sQ6ZtGSNJtRUF8A4yUnUqUVpnnYw2afHPGxJdp7qrlS3LkIBdVi+t
DxqRdPRPJFtgpJSTJBDdzy370DZTeTTpFU37v7uuZ+WN10ib+NOwuF7/l5s7LHCJNl1K+W4f1bul
rWOqHAqaflJVlsVJJThv4HFt+mMkZ2yRuPSKzODeg10Kr5vKKFnN0Wq9NM3X3g9n9P6xg36GPYrs
N2CTSk2QFucko3S6poBn24J2XSRUZtPbfMPOnZWLbXtK3MfjK3a7xm2vM1vRzJmbnd3/sLWfJLwF
bcETnolkifgp0Q5mOokSkVFGaCzj8BQ1yLeaMK4XiGzidgIfWkYxeG2wBZL+woHQvytcu/11jEbg
g3sJKYL3HSnnTTkYWE1WgG8QK0UXEmBaJTLte1y/kzrh5VnGS6G7W+FWSn/XHNIs3BiUz8zUi0Mp
QCGK3qLQjl6ctsTBYSpPRhBLabKUEqjhe3pT1JaGELQw5XUnwh0JMwEgYFITbwYMZSKYUw0v6a04
ttnr3wGVVdTMppqDJoPThWpyLnq7oLXy8SYvscQDHIpYZw4U0KhN41MK84+HjS6AHh97gKbWHvWr
kPBMU9IeAEsmJHgmcpuHRVtxNYpk6TZXR3g01hlbCT2QGvvh7sT3vX3qmpffyvYkJWxXqdq/NB57
fTsDbmJsvs+4Pq0DzG3jK/Mg+4EXwlI57ARyAoxZZQubBu4XfXz8hPfPg1LI/lyQcDWcsMeVTvoa
SOnmuqyTOBw2lRt9RWa8+hJ7BpD8mdOxY2MdCwB08/OGYBxc0VDWc3lDia9izb3sLMiLK/tinZjm
kkKy4qUjNC4hi4wJPgCW/N2WilP599+FRGStnIj/Ipffm8cGCJ7QxDd3aY4OqwW32Tayo5IS2oY6
LutYaXo+FPsyiAFFtPr2t9PeDghedkAATF+CudkdL8c/MqfLjsszKzykMGoiHZEtKFxFPPGsp5d1
f20FqNUKEYDg/Q7WcjHZjRXd7ANdd9F1Ku2MeHxJEpNcp8Hxwa0Pwi9YpN6v4otvOK2HgtMhN/F3
vRiJnx+U7JL3nz3kj0uuBgIgRZFbPY6cPo9Umeje075MZsha1m/mF1cLNVz/FXPmTpPp06uw/e1X
rVQ+3Zc026Yhv3/gxZgQvT+cUZ8KRjEurT4X28VgtAEJ9Zh/qvDy2liBdTrmPSJLUZ9xAD29dQYO
OAtRtnJ5lYfPSPv+jj5a3MvVo5jL6ebKjY5Bp0wr5GViZxC8jUhsp/HBtlfbflXbsBZ0lOkZXghV
bn5jOT6CR87SmHZzDVC7wXQYhWG5HsiYhXumJ6WHt7N64X/jhss2kiUCGuzCiajqxHiISd7b3l4K
wN97hV9MHNw6Ojbyrm4KYg9YZQLLQDyi2UFFkdY2jnCXqg8hsSOIF8Q0no55ZCrt9CFAV2QCe/+q
069L8HyX4SW4Dl5E4nARp1/6fXmsmXXzS2Ybifye9iTkMNTOYzaZt9HTXG/VlxnaK6J9wV20RAyH
kM/joae3LQW8YV0emvGeZ+hfWM0FCYgCyD8zYpiwp2XBd3+h1yDYtPLklElaXa38MosopxY6/OY3
Tm/t8r/mB8GR93tlDUhqQnEPK2a/DUi0U67bMcVWr4dJ+2z2IdgFQMIunBDsqyQ9OJH2XF8QWo8u
57UOsX/gh1FrECojivLyvX1dsAt74aIaLiTJ7QSI0J6HZDyBRnI8662y9mU8ocnyRbd6qvi/PXH/
9oFeoHZMrfZsyo2Z8Uz/iWRSzJfGXa/S20QMAOy2G6o3CxOSPTpKgjA3EHT+bZRMycDDxGMmkeTG
4nasWNzvngRh/kmGJSpi73/s8GpZrGv7TtbyYObr/cd0yUE0345lVA2sR5HUHk4UWwmotZWfGwje
BuyIRDEDZ05isO9Rt62xEG8tSRxGSp+/HHtU4rUEECQNAXWfepHPQZxQXrtWXsC7bUYJzAayhq9f
H6oVTYRGXBFEHCOGWq02qQ1V6EgIrxukdjyJg7+oSNYQH2gO09kJRx055RlCrr1MllRsEEWuKd0Z
roWDw570lxmtj8McBumiMLgPER3BzcdHw2SDu7rPUuqAgG6sdh+XXQPFf++34YB7k3yGt1EevmOA
0QAlN4Ze8Zi6pG0Xop+MBNKCvsZIqJ22jLEfVB8Mrp/h2gX2DP4AMewazV8OxvWv43af8oVHoiWA
MNVFZUx++AyruWt+uDTFwBtm4PvzqibfbfJ9nveWjxDb0ESectNcftCKOQmbRptTkfZD4B1WGVzU
Ql/3oXgQre5P9fD18TH+Eq1KWWQBty4dNxABT8jwpeqONk+shEqtNpchYqIQuR0eababf03JIwHS
42MNa8yLDbnh4E2ofcw0huyW0vuUFul4FmTawUXQnebrUlu2fsobkPy8aDTMCdUmzuXTAdesGIwT
bYwrIBb9Buh2t4/+pRPaRFLIMpl9RGgv9LiOZCQ953PbCr68mLiygYjHVVwnEmvs5QtLEfaxp6sW
wTumH8mwoggaaN1Y1JBhTEa3UNZnTfF3heDhrabSSsNh/ekSkvUdGG7/OaUqFcXPaXSghKhvNAnT
ZKNgZgZZZL9UijtBAhQp6d3HQ2gYMr5HKxBeZEwg9H9+RiPhPESrP5l1baC2iRjtU7hlHnW5sKG0
VypGOcU9grV/vYZljYgrV1LYWWYZPT+uC5JMtUZufYFSwEm8S7Z2aE8GOJWpjwIQrQVuAA9w17SX
uYZ/Gn+/IMsJ3/bPOpj1PnxusWePxLlbw61Nl2q5zv4uOAz28/6akXDR8La+Z/9Hvce21vFqLG/m
ZmxTVpHVvBrSmDQYt7nZMOj18p3HQM2nHXF7TfbdwiUBN6dcPUdYhMrPsPG/RXSmKM5k2aLWsTNV
BYpnwBZ/6HnKdL/6TMjkdXZcwpz51d8Z0K/q2RSGaskRsqfgGspg8m5ik4QG1RUJqDIyyZT1HY4E
hoMa7Qg6YeQ4/Ao0oyuzgGfmoqIIpXeqFQEVvWnHT5BDQgYFa2C1TO+aEs/7DIN+wJb9+YtRDNUc
VsU1mDRVMCai7kSExwFWfpAo1c4mYwlH4GAPITWjhOtwwD4bXyQE4Apf6bRTriL19Sy6/nH8q2Zt
xlNimW+DXW4dhjce6QEjDVoggvq/IbySoTcpTlK/k6ePlfsW6ht/D4fPYAbblt8ZFAZiBWsjIlRp
mvGKvfZPewW5WAY2md7caL1oRi2hGDbbGx/1WfiPGZ9TbMxGrRKOKLaagssctMFcwktQck0UA6Kv
aMH89AkaegjqwX1JHWC6DHV2B41x9si6ym6sNdc40w5YsxAH1rGoNKxsqJhq78RA1t/UvQ2Cew8n
LmQudbfFm48uRp6ivjfVcvMM5nWtPpQgmQPE9SgU5X04aA/9jJHWHqkEs4jBlSZFK5OJ+c6zwyC5
u+OiAua2DT3H//cfM2lmtPIYrefihm1d+WV6SqT06BQoI0Diy8u1+Yby1/n63u+Aze2vwo5SRU/z
xMw3oDBT+qHYrXLz2piL5NOpPasK8L2nnj+Xu4lD0hY0UUEccQjcOrUdjpJgDj13XgNU3qzwxfWt
UZwciZxvgYc537NudP0k50TC2hX7Fuy2rrEUcZbjbBQgBId7xSY3q6esh9RE6q1gJGrspSQi5/E/
cTBHesdgH8tcWaIC1UzgAX5FjymUCEHasEmxDn4s0cXorq8mjkIQl6moIUoVCDbeFSYo5VNhkhKU
3wri/oR304m+mueHbJ/zI/YJjBLx9H1Loc/arRRt7vBUfV+hfZ067FDyFfr60lNElg/uCGg0K88q
/ALhOvKA5dVNI5ga2RovSmo1sqn1HI6vaHfveohoG0MGkK601UtXDHLI424DUKTlhemns1LiGs+p
lZP0cVhiRw25TV1RONVsEHXVbCiT6PxaGkO7rc7u9bohcdXiKFVFn7RKkQ/daTAJlN2UvB2AT4UK
E2l0ks4QPBfJE/JQJ/j1XDCrvuHMtwFSoOzTVJI7MNEyMyEFPbTs4EAqJfH8kbvtnb6l4rWz90ZL
wXgwxV2mR3G93pm/wsElpRzjHwHCiwlxZWRLGMLVfcYUQPWoh2P7m/ei8IK/e3Vapc454bF8xNWb
YPSv1XXvx/K0HC1IDGw+ViMoM/gT7yr36T1k5ao4MUdmJ6XjiLbjJZcri24wOXKMclLBbDGmzw2H
cVqSVIlRHTOKZJV93C8thmgPUMhLKulbGI3d1KrrKYgSBOuvV/rymGHDiKxNRTxVaiipvW2iK1IT
NQlPPzw93WClOqmXPI4v/5yWnTQnx99ELXCgWYLsX6nbVJii+sNRpQblEGfZdlpo5FKbgPNYb1ac
u7BxKXA70EHbl9UpaoJ2OhUzfVZdvDryxfepiXFK/pf0CyL/bgwX6pu59H8l57SvopPHJVf9qyIV
zQgOq6BfmSLe5axBhi8fV4HGc1zixI/xG76IakTIrwJkNswljnG5iF0/t6JdfuQ0VaZXjDT3IQwr
lVy/jGqucJw9pir9Qxz9mKCufINp5xzrcwR1d10zhoEbsIZTsBHFT5PZvIlXdcGdoTkp+2ThxyUc
4D2cAe6aCsAZ74meZ3SNL6lmpb97cHDOHyh0gMzsiFESkBex2rtmbhh2ydqz7Zf2IT4Q2XX+ZUMt
CHuhaalsmdDQw2q5he/i7HjYD21H6BxTGqsuE9sYu4AGR1Z/hrGNcCjYRUPWyJirgikpwjMGgC6e
pKTcpBEmr78iYtfLEo4PwDBoCEzrnF1oexbSaOGQhZhhRupSsL1QqEWTfc5Xnxzu2L2N5TX/Sylh
kkohmCHbOZFXPs723vSPIHJ3x2p5HwfF+czhwNDtEMJRLlegsClV+7SWuh3U9DZiY7pnOpUz+2tm
NkEAum/PdojGJ+lXkvRfv1x/rEdGgy/JI8ZIzfrvfSd6zLRKVr1X3C/YnIRSbisVQWp917hfS3dM
gMQ0WZzXlufHRU68svUQdxCl2KBNFb4yFu61X9xdrM1Y0efunVqg33sYlOReD+nllkhfBJRfhD/r
/CiWbyic5D6E2cNo1U6iFeJOSDgND9Xp7scuXP3WZo645VVF6lINIY8Z2lemXB96wj3Su+6LtDZO
VqPa2GzS124z5TAzPI8AUxFfHXMirRIUabIhsjx6hhGB+H4TFFjao+NnkgETNxVr8pzZdMoevAJy
6QqHwaZT8MZHQnI0KnrCqtApIjqw1cJ315jL44x7JuC5wTl+Bsy8EQ9RdK034kLvCkzWyDcf4Kly
d0J4Zbi1SUdhDR51wGJpKAhiu4aXgTrFACr8mrmbaVFsIXvnv9l0u5Dko5y+tJ0BDgL9Jhu6KSwc
vBnuouMWEEqWxVAHHY+YvNNMIQ8qmotS1RnaFc3Pf+YiaQicQsTrMKfnCDW5uLVcZ896LmO0SH83
cV2sfMbd2QWgoJn/ucdh6y3GNz0VkqrwmCpSopiGtCaJXeJZQ3DTrVw+M3ssP5Nv6AprEilW7J9B
tZcbAANVvS3i16kbHZeRU5nj44BOODgq4bxuWnDRCZqYZ312qINqAuD4g65fD/VEvif7c1H5TaWV
364StkNC7hiH88a96LnO41qGfWCfVLRpK50+UVFFIpFfMCaDj8Xx6lNgJ+MgY+9golHM3pcPT1E7
tlg4tMa5bB1038DaUBoMu3KgQ1ME+P6rqRKaiENYoTWIaKG8wc7Hs+Ng6Ymarfh5Yift7ZY402Lz
Lg0+XviQnI4Bq9DPwXHfNmpZ45os7gMbuK5KOoEPB8hsdRZPrALvt4F/BxVsBozjOrB0fR+GyePK
8qQB3pvfyyiy5AK2iJR50JtLDAVzBFuolpTD23FkkAh2/FP3Mu9KWAVjqiulaf/KCZXuzvxtoOXL
8rI1xr/jWgW2zvxGxEy3geqn1fSk1SZ9c5Wu86PGczzaQOfgAmBPZ87CHcNiOehoSO4MNWmZ4ACU
+KqKWmkQAs4+OYTQP7bV9Oe1194mpHCs6Ymt3qknzOf9JLgHEFg6iPqBmVaXU0jRkhZ2JzH91bQ7
kgzYZ926oH4zW7+HiWIjyUJF61JirwZr3FQq0W6/whWZ+uGOCg0m6ZUQW/qMKV1ss0cQQq1+AStu
NFhq6yQdm8mSGfl/StVvmpX7qoAN8stniqTRK0MUnMtcp53d8doQBYhmND7k74taongDYNVUtJSd
obnEl5lURncHOsJ6RZeoxDaYM0uWIKml4hsGdBTtBK2z6VhQx8lZwHLE2M/OyjU5IU5rRhtMjPlU
92DPkem1bMWZ6hL3cxOZVu9TTG1QTMWaD+p1aT6N6RMVVZ2A27a/mhQoAaPDhBomIr44e0NTutpK
+ccpdheFdSZFcoxiLQAENFbhcnwp2knzE4+Ienw45OBgafbk2jqXsfefn4ovGfcMsOvMGVzLXrXn
jlYkIPs3aL7NtFLvtmoCxT4ZGWRj0w3P9BEJhDVDJ+9qDyZwtKnA8JvPSq3/XD9FDJpBwUb6KZJS
Jq73UUtx29J2frKL6hl3CX8rRIKK9ALP86ftufuWdm8P+cWL77HJctqSBeabNC6+BRerzY0vDnmA
jIFFzpzJjZLaffIZJCCqUo16v1M3cNsCoBt5CrTy+5pSukRtWJqKbd8mBbDyIRVX5iZiH3sOyMj+
ZSgrPBiC+o8lVUT1Opl8ULYbMsjf83+R7XKhD7hfIHbocvusEfHg+pt45byrRjWaIhvu7PkzKDdg
1hTRT1+n5xpvbtNQGSAvynQD9ipIJ4iC4fBLTUmp3ha6Xj0B6qmxUF4cr1g0RxoaescFMKpKOOta
bTbkjA4JoivIhnzRk4TnKJhZbcHRkq9cBpAibnZs//P815NgqrzcmII+LgbdGYkK9DErpEbnfRX8
hPfaktW2S9X4iRwMl9bmhigs/ySakJiu6XgTMJpMcUwpJNjxJqVf2g36g1Z1f55nmLp6z3boKMLQ
ou4KP7SToo1Ce3h5sALDEXUKGvkJsdDKpZtNOp7C6kRfSQOyIoY4lqOv6mVi6n5DMJBCKY9xPDD/
Ad9fqixHniMSAJE02kzjiml9jtkLv3LIngZo7t8B0eqYNNPT2CjnDMvUe8BfoSPkiQC0ubgyTRVP
A7/wSTpa9BEB6bdBiQjOVEGBrrZZRSdtryurGFbgs7zNOJnk5WInm5KLLSCfIgy99CPIwT5p81BE
9q7ooOrgim2gqNZUBqaRN2PoTAHeS5vJz7OGMOaJadAvm3GfRnyuoEC9qa8QmirRO3hKwoTWe17V
3ENtfEVIFr63jp2xEh6/cn+i+K+T1Lk0PA7AdO2jdRIAufhmHeeZUvt5/AlgqVB2q5E9cspn6OUO
MXtzFeu2jFDX2KdA7p35DmrOKPrdVcdt6yk3q1uAx6lqkX1oZ3476tc0SRfw8ay1+54H1JdrOgBG
3JSQIgqqTuda5hTBavERWT4gEvBOko7mFkAF57zbq4AzMY3jtmfaBD8SEHARVKY8GcWMAjPwB1a6
eLwBHJ3fjh1pdFZ/HLZSNwQw+gMvBekO4f4NbYsb3qh80G1bbQHikwRLQbhD1RVR4GFCS/Ab9Uf1
VUIfb6wGSx25a0j8Ngnkb/JhpSGZ48yLA3WvXPxJALfdEH25ta6KRjRj5aNY9mpkQxxNlX3JYM6N
N9rKJYnlRufRKUidrQSR0uHppTSyhXgU4ZPCEvdcxxFWosvXl8id+srb9Pu/llXimomrlb+OHS1E
csHO4mwiG+zDLsdQoCNXM/IfkhO4zY4t3OH4TgOR86mYt05py+fStf+rlZ8wjrAY0Ndt5HqXR0RR
xT+zta9i3COZUS23xt3URlPT2fBMzFMIXr5aQx2H9fJW6HyLIYNPyR3H6d59zzrpfenD1KK+j7c5
2cW3sFu0q4SeDtphLxmsCpqg7lmdMylhlu1YPXzD6runJexpNYSwFrZOPDiabcy577DBB+eVE7/N
omAsUgb7K32QyYumS4JT8un9X0EzhMTdNkreV07zNHeHTy6hJAjEl50JDHRAw/yjtxGvxW79Dj62
wBQ0JA9d+lqvuCxdpk4FdJAhstC4xCFkNsyXrNdPgYreVOE+RVwztxv9rnAmVP3TWZ2BQlbEGJtw
8e7iqvW/Dzb8I2By7zLSRWKwa3YRCclcWqBDq+kj7lLk+V+0E3TWr27F5V8yR+YERepf9YDx/gMh
v9D1V9BLQeVoUayamXFGCsUvzZY9QxrJxFqqvlSQBjUU99NpX4NB6B4MXTdP6gt6UmtBfjyKt9JQ
ei36kpfxYOpWCgazfP7nYXaCEPFGS1M3IcMt+nmOptW2MhpNUBYn4SGg17xJOf8rpf6pzVDSvm/J
rLievjuIUoOGpfj4fhrdbnQvZir80M/UiCYK5/3RRTAiReaWNLg2sznwGeCZtpVafKNRxwyFk6ej
dPXe4W3qsKWxhy3rfYxxOvmYU1OOXDn229Ka4Kqd3l3HTfGpN90bk8IZXKy7wZGnDL9kVZVAvMUb
1iXJM5mncKc9SZ9OL2hfuEctDVy0FIgWYYVEAszmMh0g8U3txo31RMV9wYMSlPXoR2f4Ef2n8gkC
4fSqhtz8q8Gbid70NMm7ykuVZ2JO8kdeYe9AVWZs/3m0wEJZ4LbVSokFD2EqWrmwi2TdPS5ioZL9
ZLHWRkbDODRbPeCAeUpNOQT7GLJ9abT4mf29HZ1CmRZuTGjZ5FqWCvpBQCFhgiHyv22xhMxmz1Cu
StCvUjKE38kvHQBeV6mCcK/wwXQLkrndz271NEAKdIcx63f/P/7V6YWlf5MM0ocEoxpwyye8m8Eo
E202EbGlaAMM994B+MLGttthj/HG5XPwcpXalc6bbYAK5bH2WcCDOVrgg8IiN/fTntT+IkjtVPO5
lsYYYN6LMCX9erp8Op2dkjRc/Yiu0I0yqU9wgYQ036Re8GZj4MJeF/BTOe9KVevYd6WwtwvqS1gi
40MoNT5WmDXxM/z9dgshnEnPZ1ttRCshMttj/9Wi0YMFtqTb+qzLQkecnvKYyNK+YWaLdgVx+rGE
EVFS4DUYQNOICsLHgpKcJ8Nn8oR7T2mLtjCGSZDpWpMCouMZJEXVaUCaCY9kDMXEUFk+XErYkQ1V
e4hREww5+XiUSKuxFb4xrYnt2p0BvKPS72D7J9eIgwFyQTh34v8idphUjCh5ojOHXvWtdF/DZwuM
cbG+oXnYc7zl+uOKtQsAJAPXUBOG2S4IoIWK8cNPSeiUiULrQCl4iWpiGBhjblTO6Fw9L9QHpcU8
4XQeWbc7i5IU4M5b9vmZ36YHW7Ee0Bupqr4MQYGluSGxryzjubRQ+vpqe5Kafel0qrdq1+U9aaL/
FGBQN3CaWYzVXu60YHNtcjdHlQwDUcgUvQOcWuUNwvqTIaiUnc7VwZ6kXSzFkEuymi9pUsV3fvky
rlM8Ei0jBPz9YqTGEt3W56Vwo0UXREGFpsjOiFDMDzL0tL8NARSBV37KRxkI603wo2hhpIOcXoIB
zGPzeAYV6bu/doJP5A11EvgI6TvlVA+4EP7OXM5Mvtyiyg4d2P8r9f/e8NuPXWbUmhrwjfr4tUZs
ZM8qgm6jfNtuNL2c/opPljqfuLSFhqNJf8rJRionuzfHVG/+IKr0qDhjaZYNkks5ryUz8B9/pRRg
pBWfSABIUiPB/ZCxwFnKagiA2QLd/w6sdXFt+c2QBMQ0XihZjpehujydsjVTXFJ//lPFMspMo6xH
DrYVlXqa+Z9y03fViakd8TS5AoH7MJuTKjRO4WscfaLCtucoeMuFcIvkrP1x+FqwUVgFx65uFtdV
kBdrDdZHHZyqg/c6jdanCT6pb0UgSfGwsI7OIEykvGpQXkfMEL+zavGKo1QKItn01lmDvWNwlUT6
pEB0MlB7SH7Jy3gZajV9ECtyu6qFpLDiAICyHk1aKFBtpPjoAPm3yTUIr5C5NVhSw5Pkx0vre5jo
qgnQGqZVsihbRImrQJAQY+BRJcM0a6hbg8wIP7s/2zuc5qMCjUzZkWKCeUC83wdcfliH1Mgbzyjd
PHSIWqe5BGjkZyuSdKZgHCLytWX0gemmKYCrQy81seAwM5FOVjLWzYJ76+RNzyjwDz9jQ6wxfZqg
FNXOyYEcFnGbNpAUnVwANWQdql3NLIZxLHmOXs0PK93eKPHnu+vK8EeMEHXuSJ5SCPspGjmgdUWH
CF0/XPo8sJo2vs7r/88LuLmkShdES913gTsfYsjY2E6Hn1oU1FhFp4EMMbbguTxyBSdj/6NHKID0
S7NEW2a2dgV0h6irfVtog8oIeyVWAhsGSWQ/v/urB/d4p+Vd5gZFFyZwJxdqCcWxeEgJpIcpVYg4
nsEwDCAhZpNXoj4UIep75S7XOHrNCXoUedwcVvNKVTkNA9Ab/U8BeZtPJ8Oefy1ZugigaRyV8epF
0q0MdysZ1jg+eQXQOMACJQn1ODk0uiEopur8lJ/MaaqXxOBWFCsvx3M9KOqO5dEHFBmJ7KdajgKr
gFMHZwXAJzYvcM91VxpBG3cPHQDpdUwlhb3+mlsuJ6evCKfSdrOViztzn2jEOxIKaL9+SkUhXbrE
sWSFlwg5XxMnpH0dWWIv0Se1uJGeeuL7Lq1EPrRSll2gmFkRQjoIg8J68n2gXdUtuurNvd1E4WTg
LrUq2Je6ncEK8fqnuO1h3XaCpZfn3h8f5zvStd0P1aNb1drc7SphNDE/RahacOv6BeKMk45tNYEE
tYVehzh4DQzfH/w9Cx2+6gAHcSOxFFoGywuFObehYA3gsOdMDT1oRO6cJgOtFDADe4PuDBZRIRFP
bsBN1ETNfDPgUO7kCJRA61vlKvuj33jQoqZxHMx8miZCLmSdBibVbD4VtNff+Pso0EsGv7hMW+O4
JSCVhpKy0zyb0/tVxhvw0fsvevorKDuinoILG6PJV4leR0TZCZXpv3TBjkSISc5awaCoPNO4k/aW
ezSlYPQgiGQ7cCSMwOWenFKxxb+V5+qi3RZ52x6irsia7ilLAWMGolJjhi4LdQG+o0Z2HpO4es+H
tPqq4CfQM/I1SPfG1rBIFtRkyQn7HOc0pkLW5sC1567+sq2c6SmaMiChV0Fqd6TSj/HfReApBUe6
mIg8YjPCW/kRAkqhvm0EzA0OFPuB0pZT8H1r6yRgKdZRoac0Xr+e+n1LAqDkYcwts+pYEZoyKVc8
v5KucywAdUoqtxiMAfkn9TE8jQFK5R75rgk5W3N0OcxYHkezYReaiZLe7CXs4AHFersFlp2/293s
HhbfuGbhhGwTuC3hLPmYYeqs415CWdIH/7g+HdkZ9gjfSXcV8sGXc453fnX08AvwACxWagOiA3VX
mIFj/qJ+inJay5ZLkE9S28+t2wj6YUfUmpFqLj0weJEFQRxapSUist4tG/vTMONHDpj3sDVP8Iqn
MYSi3wkDgrbfIEPWzTSFHMr2dDJ53bg4oVTVzkFkYc/Y2soIRuJocoD6L65hsl4H7npyGNkMD/vl
Y+xJJSZQeZDSmhk+KoBA7QHi9IqRnOkUVLSUwrATMEJtdAp8eCVFNVzUA873v+/X0agm4dE7l2Xk
RXvuUryJYiJgaNv+lx6IQZ+ZJn8IN9isq202W31dVKcTp+6Ocs2swqftI93v3r9mJOCOXWtZyERS
098HQT5eFLtB8/gwxkLxGn7trLPoawRTHWFfOIz9jtRN3fVBQ5i6Eu2QcVZSMYdMTxXdj2Jqedri
rYZNymkdGGkBGYiTXmBrWuygiZrYaNHFAUB1V4XmQQ5RbDpxR0IP9FbQVrNrI2rYE7BH9B1Zvimg
ETFvDN2bDpTNFFokU09iGlcYuuCIcKCjvzz1g+QWz1+x/bcIkvQxY3pC1++LQruSxqhOus1Xg62P
UC+L6kBZ4/4cO/Dm/Uy3BMblsMyOgMwCpTid12pCc4nxePqgrYmQvY48s0BPCr4E3htcFMqigO9M
Thaybt1bv5DvnHF0lmkZ3jLrLCQbOC91Ygu/Pu0INgg/1YLeOrcCxSOdujdtJCMQznEFWQV41ROo
JFX4vmmCJ6rgXVRJVlsszQhVl7o67CE4ApRMLdjaTB/8DeNphZ5R3drbYY6AHbODtjjXce/HSE8u
83h1L6qT5goHUHMjm1wn+oqA1HGGLcBMzGPDa6lyDbxv1Q1fXHaztsh4xODL6/oVQVupX5IhlYo5
ff4J/V1chuepLEv0XqJa8jT63DcZOd03AV/v+wFwWDo3u3pTdlAc/pBF4/vEf+CnjvAZR/TsgRPz
hEoaYK4PGYHuUb096qP3aKxIM/TE9mzLqLlP0MrzqeeeMki5iX15HYCnZc2aMpW6w4Pe49AnNws7
YSHKEPMcfr7DncuebdioHN4hesj03p31iMab4X5KhW1NVzYfOqE9Yf8smzBSWmXU2tZsUF9GQPLg
Y0pQXF2RMXXSXQTSuKSu+O3rTaXmaHCtnVViMlMs5qqJIPif9spMl5j1X8JqvNsn+Jc1HERj4rsO
rKqiMZGvAy60rxtb73nC+w8T6w8JvGW2rysxdzey4IDtBttCiG7vZvfk6tT1zwvPnIKweQghpQaT
6nnxx502xzSe//fqh/ZkCaOFwWixoh3P3wpogB3O7D0OLE85FH7JXck3EiR6PAQPc6VbnJ5qWg8L
jK9UkZpl1KwsZylAN5Cs9/8MLzOIhdQbJgmj9j3ib5akS7HmJve2/upuqNVeQq+or2sOKHfRzkS/
f8OFCPA1l4ywPmOpfumsk9Zb9gnTn6Oa69e77mPS2XDYwNvDD6JXXThJkk3evocr38yD0DyJcSLZ
emYMywOAjclfcx+O2Y0O72qi0UMVSIYxF/oTMGztWff8WjxR15Q21b7Vn/mn3jT3XcwxFMN+IZOc
WR98xKYJn8+0nMT2mr1RKTMsdMBS+bCGj8t0Ln1x6YG3fmZZcCp0QbIpcGMRkUPnhNav5sbIFUoj
VajfUC+W24kBfnr/iizjHm4I8Z93gt4JwLSR02C+x7eqDi4mJxSVXHg13T+wNfmJUNOTfzugQLXn
HpAZgA0KgjP2zudJhr8X3Zy0Ij59fBqMdaPk0uAYX2ZOeyLTEvVl6rdKhiLgAZxdCHTyLUBcpRM/
oray1fycbBbtzf+mY5vgqs9wK8rdKz1jUtTGoySjt8i/k7YooSattHzwCIi4frBcOJTpg353H50B
FuyDzVov6Zaf/F2o8X/doujhobMX8U9T8lcBxiZb4CjjHzpM2UPlT3uLWksATxPGMaWChPXrPKoo
FNaVhA6aD3b7q+5Lkk/hTqu7vUKCZSPwL/t/n1uBc5Ojnqw+xsorbtyjHhTm9BEnaQ+gii8UCDrY
fe+48S1MVOhkuFiGZFu7SjNtUdHHbm/A/0b41nXc5Jv2xtATwvKzweOXwB4sl4tLQC0pCMfQrDIs
I+5e0YYxl0FuNhbe3/Uvt+K8rSdDPGnCMXY4fXvpk3Fu5EJAwm47nvwyBVSmhTN6u92pmAw2yhIn
8wRdMjOYobjZnzB4k02NvR5RI26BzzFBb8CHIHUhHJc+3TVu5xVMEx+Kg9MuPIZD1zJkJp3L9hw8
nASZlapy9M3+ShMxf/byMRHYNGCx0yqNhiDeQUI7g6YtsIuzffpJG5x7nxsLvXCKMUKCGJa0tyM6
20pNzUajyo8KqweuhTHMUVyhObZ2vG358ng5EoO5NDM1Sw/J0aW94MrY6s/fTH3UsvkyJAQeZuE4
1Du4GoTKn+eo7B9JKMbvmmei+wgsfuDRpXrYvzblGUNe78ah1VSCsaEqhg5BcKueI5BLAKBtRTMR
6RgZBrLGknkCyuHprtT1KnKmgadjlBX+ikbtXF9K7nU6B3OjlI9NmVzBTIvBiyNdepctcXBZYFDp
Gfey3Mw89Ea7rds6pc9CsF10HvNTvnytQwZsw5kvGzQzD/W9opHjY3LYka5CTtECJf/gIdQcQPzq
TfEKOazEm580GI4injNf+Z1rCZ5pu3AYKRm9KtL48yiE5JCwbnQcaTx0/pCsf6h8ZbhqWDQ/yvMu
r4VvzDwGxIQL/SNAxg1o7A5nm7P7z/PT7uY1P/t0MU5mK+arYFRdtc3M0pCSoev4KGF6iihkBayK
6qnQTo/pgiUlDhNfcCb0qjM1X8cEDdz83ZJcUlGMnt/S95vt0wxoAnixI8T2LuxqkC/DrA3ZvW+8
12vqz3Y2Zw75n1p4pzOAomByJDhgcJF8e9+hyGiIToe7lzVZzzUPFXcqSu0LIHt4ui9aWC+SKHYj
o7N9J6EpJC2dmv6yXu4bjvu5tgWCGzr1mpKbSwIKuT5SWT0Iin7BNZKLDqOdKsaX3uVRBp8EcxXe
nYfLdnFup0gfynOwFwtlHLS9WkHJ8FrHCWd07K4SrdfH9guqoyVvz8+02qqGteADYjnWlU1EdJkI
/HJai4ur48Q28TG1ge3F9soOq9uHqyr/+D5E/aU08kJkIOPT1as/L9AqMCpySYqPRu4k37ZkAi5P
MQMM4HrK451Izil5Vw5w9J8jYutvhwFzfvpslGULW4tcHNO+jIPcipGZgenCkxyCDURsxUgBzUzZ
tBSJ2399k9clkd+dcBnNM4p5m1MpMYZuRQ6OGhUU6VyyUnK+fuV6ghQAQUtr5oV2PxsOxdrAR7js
x5TAa1ihcxTja3ERogCIxSiGpkf350GtZ5VvETXGpg7MpxMIVwI9zJczqEHGT0cpOn1xW/iTUQbL
GaL2/lnxBFImRQItfZgsieESPN2SMtkQQiW84i9XsYonhzlYZZ21NuihDxYlftre92zEaw9G7MpC
f+atD5W/RG0zKPUilE5uxbVCDOdjJ7qc1ZISEJji0vbKXJ99FBaRwGVwRKug4llSNJXcOv42ofSN
WvX9io+mq4hkiKqtaGy8yQNYiW+CmGSDuD5mtDJP96VQJsjK+79Igm62z1VpjtG6uXRitPEiJvlk
fbQ4JMaERsCWn7y8C+Ei9WIpv22Acn6rWXeimX0z/Q45pGxQGSUP1eBOZ6om0JQVToFuRXJHElnM
Zcd1S/OqMHnnbmNZZhwphuvVWCnEi/BqRBnGqTEFLjGOVvt8U70lzUoMf0Va6N7LyvXpl4HvbKzy
tXCRAkT0Nvl9mhirG7ehaRopGR+X7cojEjGk6rvsEHqvqABINmmwsPSzd6pQt+x3npBelJBC2Hpx
ez7XITShuYtm0c33gGL+NC3hv8T/boGAIJHs61nbNhSkopEn3anuXvlyJFZjnWNn+ylzyHxpcIIR
6/T5KtGcvYW7P6yi6/Rtte1KISjB39JKb7cEaXbFQzRVJ30PB4gx7BQ0Caw5gLPRU/U1dchFTxrm
uqsX8ZEFkxxGGfIW7KdjmGvAqq+3hKD5tV+ebuOmY4OKqc6mtk12XC/67uO2lZ+wdbaWYk5wU2WV
ZDiUB0l/RIYdwqfvqx4oNFNTiuxNhfI59cN1n6s3yvCmVvc2LAMCw7kCytOZhRGD6VyiKOz4MHRP
Sk5LDboa1c/Ymm/Z9oPlqDvlvxDEcGyWpmwx4B5dHqGUpanpOMejwcZ+bDqnX/aEHF/QXg36bYAA
jl2Xlk9lbwd52OiviPWPZVOtYQWi2jaJZP/rSK2jRsbsgEvz5liiftrZLvhP9QwH86RPQg+asWo5
mbtAW2S0ng2jCncv1x/IXhxRTPHPGSYmLhOshIklBi2/QR8CL5K5OzMU+5JNLmyclYHXi8eF12Ee
J9SCgrSmomzP9m6q5tOJSsbo9nAK3Scp2SjyYQLA3eW6WsWdNmtC51ncgX72tnGK3JHLz41KxhDv
jTmP72g7ExvMmDyHJfPBBhDb2Qgea4qOR8YGF0Sl9YfAk1D6X09hboBly2rgQOu/P7tRkkNim+p5
x8CypQlmO/Tf7xkSS7TiQI7M7NcyXQLnxT4J20DXHD3ZXfYfQlnKTvFiI1RQOLmtM5t8qBnGSkVl
4PClHVFYM6dDhyChC9QEsrYUajLncXneKHubS2wdlFIKMFiOXzZWHrtLw4Ing7f/y/BkL6vdlT7S
96nWofc8hL498vkEtysrvOAdC54/pfDTFGhYhfJmQ9Mt+yUrLTPd+fB8mA7o+cR6CfZSqpZpezUk
w7stX5+8VVEsel2/75H4Ez7zLlEGxfJFodPjgIZSNLyOLKNUCxRnTFeTmlbP2bjW9qZDr+jxal84
/kdC1kL/vSzG4WnWZ3CS//mkYpqfZUWuM6uE1PpSHi8O5TVRqYEfqdlB8N1apeu5aMG1Ng3NgleS
OYbyMTE83vUkj+rDm5Zgwo6vGBhtFGK/mtz2TSuf+1Klr0kRUAaI8by2x1S+kvMWEwyc65c2Q4Ce
t4rNgTE1G8D28jROt291airYI0fCZiWk6Fw97trDvcoPWvreWuKd+sUoUhwlQpCFOmUShH2eCYDW
XdTLZcEkEmOESF0RNLcebB1pkgCtYn+/9oUXcR+I/D3/UhilLiDlp4+U1j09JNQWoS65D0XI4LBu
BVx9i01/HsZ2RXgvmWSCNHofSA0JMNQJ+IorX82LhyXz05hKZX288V9rCz63J80uXNsjXy8phdlT
QISh4Ygb9RCfYqcDELbecjdkVDDuOvG/sVaABr3UOa3Ws5pKdFvJADU/fdHK1byUlClzDfB8nGP4
MK1nghLvNQ2v1abTXFaxJMCc0VAjyDXjWd+wOX62C4LrOxyvcGx90/RfBoc3Ck1sZotuPu/VPaA+
CquIQOWeCDOKtgnJusaOJl7d49oN/cramfbMbTjV+9dghUZfiueLaluL7wia+lWRoySJ3oja7jY2
TDaA3mNt6MX/X7krKv86lgDav4CbiaHs6qv50xhw3jXDqGQm++MdMj1XSr2cCqlaWRBZzpBIXKq3
zsBpyDub1/zF2RrgOQR+Cej0/cyui1qHGJT5d8x14wW+rLiVGCpVbyIke4YoKeLyFHP+/OgxMaSC
l51SqBSTcTWj4CZ0YjEUwvWQQVLw2QZNeGkmelIqPT4gAlXHOLZWW9H8GRudjgNmUs5QKHFDJ3Wj
xqLxrkzRkel24HkyOI5MquEeGK+VbpB9oMoIvkq02Yp6PlUyj6108L5zLyjmWP5XzJzYYgYIINW/
n7w3q3m71qW7OGDGQx5fV1GwY731bcceEG8O7gIraXJ1dBrzcHucx/juRgLeZY3+G52EDhqpoLvp
aae0HyEHuAkNhhWZT4jepv9jI9NOeLmcc+QnYkju4n2Q2a+6uQGpCnF93dOriAYwiDpzXJ8VaFfK
CLpwTmkCRdFQqhuz3ti3BxZPkTl0ABu/YwyaskB56ZFnxcGFo2xbKkQevfeWTdpWdnbR0E9zARbr
6ovOhWLAEMN8HLMRLlQRrHoyzCFSwRLsWyxOtm2UEsopSqluWB3NJbpQVGFJvw5r8EbKXax+48QT
E3xSOHhTmpnWaVQhfZXPpP5LnfhsXXsPB5h8a/jcf3dsa3SJIHlcp2GTS7YzfFXOGDmAaj487Bj+
zKBCk4SLtSiG6HyhLXQ5irvzt5teGLRvY9GbFqnMbYwE/WM54qZnRfFP5Rmrd6L9o+QSRuiVWA0D
W8VxW4EC1sx2XN4cr9SxdwfujdhKXd9/ZlWcM/RYOK0paidj5V0Bd71W75UGGgrjGER6fXfDn/m1
nLSnJElbo7l/V+i/8jIU9Sl8AVkrLlm/9OuI84qMpk+nGKH/Oi53mOw2I6viMQ2cgS4CZf4DgY7N
HMG9QUDTvkBGuHQXqwsNftQWwf4pTiENuJoZsh0aCCW+IlV/6AKNnWKCreAOs0vcX0oCV7FZVo5m
iFC4gac5ZPjE6GiH2WroNxrT5k1kf0t/I12hK/GIFRGyL8JHd+QlbvIJPimV1GkvTXDw7SIqONUM
iszh12clVjPKrcDKd1PLV+NONXEiLvDXkdu4ImpkVqJubwfW32249wG+rdosG3kTPsxobdrBMQWQ
xdffgyy9nC6Zo1H/nknGMRRfHkAEJ6AL+55WplPhWjZeqaBk44INnoe8+Rvgtpkmozln90BASPxK
JLkaGS9erpnHsriGG8WiL4ebZt0xEW67LBLIJKLXUcN85X9rV0f46bszzWzHASOPEs0ZLY3GBjGa
AfuzU1ofwYZhLPqGrKkBKTff7ViltsXXEMEJkLKabvtFOozMLEuQCmJBIK4MXfA853SseTO57bw9
5kqFkqFzw52NPSRBoTqYM3PeRBE3OHN/wE0aIdewEny963ujF8hdRwTJbLYeVMY0JEb8Y1iaptAr
dnrvSApu7G/aUE3eAg0gUr640RDvIA9p2a1WEwPY1MoW0oEfI6XaT9MkXruYnG2V5CcIsz7qPHB9
VTFwHVgbuywToqatvYhrIGie0tYHk8hf6Ypnsm2ysc8n8duHzqTPZgST7336GwEYE5/r5QX1y/jz
FkrsMTZzJ6nheaBUNAfps3PxjiAFOat9ljAF29FiR11O2rowJlgdcaXBoQyRqu/QqQkHmYly2D9T
0t51to7fvvr9iYXjV/OrWGFWKg1dNg73LsTqPR7v2UKpLezm5mQlIJOYXTxdPVy4dm7qRhR592lx
6UQGsqt5Z5IbgZpeR0b5ElF7YRnfiIpTywJaiaJNd2+EDjNDNKTrLOQ8vDPjmzXXCjFsLuGT77Fo
6nB8zA0ZmH5vNRbWfiUnzGYmZOuHjdm8eedR/peIK01h4wpEEtPftsMs7meaREVNsDREuPhQWBdu
eZl2v1ys4Vn3pfhQzIc/g+tC0E2OC+rHA8PHnYHNVHWbmZJSshXLbC8ba/K40/HuTPWElQTx9nyt
W3M+klvQ9uFTTy7nTi2JcSq3eBMsqZhkG+oCey/U/RQr/iOOuF9Zj196AeP/FXDgjGwTrCYzDrns
WQnLepxuldXHUngwIE4blhxjfFXKsApOtcTSsbSmPZk4z0ZqlE25tgiDm6BadwAzj83RuOxt8w+J
r5mZwmlTiHdB88OuLBnABmau6zcDUmXzQ30kzhhtF9sckx8QDWGxoNcjohNPPEHsJ+hUk7u0F76L
MOQOCNlyj57dRA5a05v0BxQvoW9syhNBoMvYzNp2apiZHarNugLlcwCsAT3uZz/hzYDP3IlBOsAf
HZds94H2B+S/VAIok90Yxs5xUQHim0X+ExidG8pHYZxRwSVQBiE3YNWTgDmQ65iq4UgjVhvau5yY
770mlBAo0TtFXLnKpVk7Q1tVLiqQ0v15ey4X09+seTEwvXT2fb4VXMA00n2uqr5PPni1du0lm0Mb
m9FbuVHN0AYbhDDk3MtSQWW4tfWG8AGjxYUP7YmGXjAyAQVMvYCkpf2106uAvTCQM5VeAklftg1v
GiZxIZA73MfUCbVLUczzl44Pu+YDXgS2X3zUAnoUQQvsE982zLBu9K3RQsF1mNHbejA1xugrhRG6
rGqvfnLC7ndMzCMIS1+oY86QSTOfh935am/c+/2/tYx79HN45dCbW0loAcUHZmCDu42M7p3CLEgg
WIQiEqvhKOpON0iQ2y923ayLPvqPP31vL8vvx8lZYPLBSWRcL/vWtoTfLsZtVyplf182eyXXAGib
w24PvBiN1ja14wh0crzs6VGcciPWNkHi/4Pa8/6B2CS/TtRT2MiOnd1ZoEEB62W2RkXTilB/7vT6
0vTd/J0TtHrAO3vm4nc1Um7uuVoBtFEK+iOy82Lr7u6eHuxXT7m453TT6Q0IjbRMGFoSzgNi6MlJ
c872m7JxvuhlU/Me+BfVKNYg9HV9KmCpBJMYBcllPavJ7S00OIOww1lv0xJKDgwLeGgLWZYKwgmZ
AYJ5LmQIWYFvfEY7w6t03b/hcm1bScGJ3+tLshXzP28rLaJz0NddiPJbFmOHIFEudRjbSjo4ue/I
PCk9BfN3uwv7HK3FvxmJ/VGaWQNMbnegusNZolCY9NU8NUIdC7goVOjg7YuAUCVwYKDQmkMqaz8q
jH714zzh9bWcz7Btp02FbITTufpzSxZmTl7h0rXux1UTqDVGjvWpvQJB5x4teU3pO2qAZY7eFiVi
IFRb5oQCb4P31rZsOR8T0POkrEha+n4mxU4OWQPCT7T8qLygteiXzDMacj/FP03aXqbBfntDuLn1
2tU38lCJdREe74ylmg3voonQ8SlCwFb9h9uEEAwwu8X87ofr9/+Bj5zpbK69T7d2dealiry3xpgB
awmkCi4UO0TVOlcMTnyt+93dYlUOUpYJAgl6pF/LJvwr2ANyb5e+csV+s0uHAo0FsezRuioEc3WF
CaP/CiRjVH4cY5bTo+q0TQgYsIkH3nDmU2+yFdfKgL5yI0lb1OIXys9IefHhiXvHVtfHQZgU2Ma3
BRlD+VgJW8VQhzrt0qUlB7HrCkjPfYHMVveQPaexQkPtNissEmlTke2wT+jR/3aCzkFg55aqzTSO
VMw01dNEKtlXWfBsH+E3FNaV5JmxJBHze+4RSqtKFvabRtA5hKfw746pU0gmjgZsX/qAReYIk1L4
OtXLAuWGKG9KZovUG7y2GoADp7BsKyA4f8YQ3574FZcZn96705z6DuHG6LEEI/IiFdEmFnFHJZus
BdYSyT3sFnBL90rZVnQvrEzW/SAyBKuLGmXqXQKlur7toQ+6vM84y8damywB546WZaMuEWxUJLgC
DZgsZgB+bRMiEBYBZjcFN4Y2DkFEv/MScJMEq6dDj2ytUj2GUi0ufo0J//gPiwWC0d9j+998TrWr
/0NcJLx8p6fcTNft5NMu6qJP/3M35duLm7ceHA8YAlOL0dOxyleGBw1BRYLYTFeBEVsuOAEaqIgy
yJAq9ozDDIGTwgrM4xa2evsQEvUhZOqf3SU4RScimFtsViViVccL6ZuYG5Z/HfojzMUhJGN1D5ic
OiQAzt+r3bsO5OdI4bGMc/b6eu5aogR2AP5aBlywVisqkGEfMLrcXAIl1QjPoVW3Lu74DDnn+tID
ql1YqOh5m9vLL2nzrQHcYq91nzhiPDxV2tKFFeg49fFpqNGjFW1d1f2pqnJ4aN6q48qO4ZnSCCNQ
iR4aQ1AtjGakRlRaia5Ie/xPsfeYy4FWRUqp7UmalSjVsrU2rldbEdIEuR19PsTQvpEAnBXC9eBo
bZXj20nxR3lIklOg6fpGBudgDuVQLru6PkiV3fClUgoF6hM+NOTLlLn/Ib/E+bH5UL08nA+1HG6E
tgjKlvT+TgvO6cambNLpdvw8JAMU8jKMZZZ6fejKdIVO8YE9BhjLJMoIRMm0csOW86tQvpFFPkcR
FZBiZa5TMPK5PgfL4xEUzaKtjb/XjYRhvRGRI8nkSdhZLI5pf+aJ5UQlxfMDq8UpzGZWz9FeLsH3
iD4wA39FpHXnoVQwxNcU2qux3nHzRQsTGeX5PNPnP+7oVFDnQsRTTbeAkGT4WQ5zp3Eyn9f/SYzi
uZx1MODXCXinp2e2hUyeMr0+ZSSBnNC4pdlgv/btJXaaCCY984HQDRkQOIgcCd6RCOEs/G2HpgrE
N8adQ8M52q7Nz04IqSij/j0YhVqGDi+uMHOrBxrRd/Tg1JLf04E3aEya0WQd8g4wGL+JKRXxMRQU
H+l6uzp7YAP0OzxXvbnePZP1L3W5NZNNjKV8BJ6VQCnBu1eoJvHVQQtGA3kww5fRUe9yVUrBW9an
62S9HISG/vSt/Hrh05xgxjIiuyRMCWhREEfv3rO4yABuj73qe4ZF4B/Qr4dicZfZkT1Kd2HZYohi
iW5sQ+SOVv6WDQ9YVYr8by1VqHgLIYdJr97/MpfTJ8V2khxpmj1MD2A8CjoBuy5BF3a6Z/w96J09
OkXjqxbvUC2nuG4oqnbNob//Re4vBDQ/FjOGkOkma1NMi/lgMILt61em2yHcEYclzfe4B9yV9iNp
owpETPxPsN1+51jeKBm1by0xR4y8xikwNKXkHp4BO+UycaQVTCOBu0eJuHKLq6FHic0Mi0e6VuaX
1D31iqpC2deTAKf3hlmdqXkpC7wDuwkkncq9E+91KO33gVNtSw7TrQZZtpQ5sO9vGaDZTTkHqphC
J98XbpcnSmRYGDtkEHMLqP1vsDO7ouJ4rx86JrVYpGB2JtGXmrFmXGstkLZY/qt6AwFRP2UqIbUG
vZ+dCTDHWK0rIP8Mdm5q6Gsys7/ENAePKHW+9aE+j0M/hu5sh3c2JN7O2qLe+2FYaaR+IVcnlR9c
tCua8zbc0Df/26D4wnasbP5Vy5U9RnxZSYbthLFXEqIA+/9PS7N40P6A5EGTyRU2BT+UmyvRoHyQ
GKcCNVUsj25y6dEn4wUvipgvDke/T+G34wGZUH682iE2kuGk97h+Vl0rKe5L7yronFimd+UP2q1q
57QY15oueK7OOPKQkLC13QIFzBwk03nx7rTKf7VOUD5Cg0iIx1DaiuWb/rZjxILQgskPM0wNVvwL
TeHcVtqkbtM6XwuJcBjMSdhPAISvpIfJ7SStG4LOlZ7uogLciQPC52NYalCMDtPpfFZjI8B7tSPS
QB+1jHB43+yR/aBV18pOyyqjj+T4c0DmNy5gu803zRMEnTajmXua40ZDd8uLHq0I1i6V3b9gbv4y
l8Fd79aw18H0JaWj2zV8c1hMj0JVeW+ued2s9I3vIQIt/xx+rnujM9F1uCSf5ZyytP4TKA2PJxNW
4jxZQoFBbKCk+yrWSjx6GiqL++QFT/LkNElhnp9oktQxdyvwMSOUHuuOEuoY73eqiyomIo8oKc3R
+L7qYOSSRUIjxgVHEfGwdpBSatT5IAQ+DFfqS6IqoMrQl/7jMfzl5ZhNbT53uJP8vMPKsps/Iuv+
GKmgV9vqFYunJuW96v4/M+exEgeUUn8jQaG9k/a9+D920d6O2TxWIcm21yWzL2+0SYsZraocPHne
OdlMj7x4fxuhm8z3eNuMIpWjKogNubqdDaVbStVy+ctl3zyGDn6L9O0Jv7yUs4CwODaEbZXX89ll
aAU498BU7ku0YUgsCObW8qRon4iKwIQHJ87F/YLOyCFlI8kC9byyhw3/Dhab3w8P+VAjQuAetXAF
dV3j1LseOvth8vcSPtTuRLSKxRlwC2TjhEnR108pDznSJC2JDQnqyPaekIo0tizb2+5hIhVwut1j
nYa0oGRtZXr7ETPSnrwplV8UlFdC0kv6TjWR7T/yyXPQ6Ajymbz3kVTyUw+4wteaPf7zdcrxj/sj
Gzqu6cK9u30SmtT4wi7LB4TiqHAobZb+QqjCL6imdlAO8qlmPD4G3/NL4CxUvE/jxtBO2vcl9MlK
9GKcKcnbyShHEKm64dJY6GzNRCpeylwNDAIQKMau+p4A5rZ930+vapgJP/+q7Ditq2aG54/71aVp
nnuE+GQPCYKjHi1NO/lZMT5I28rhXiiUMheMJql6+pLHKNXNyUhXCRxSEquk0vRI9G37deK4Lex4
8LdPo+cFDptZDovoO+s7tB15l0bIXi1t4VKZuGHP3dTuyF/XqQsdBj6p6o5ecGDcy+bx78snrNRW
DGPsU7FGuaiwIHmCTg3Hi6DzXqoOHajl2zsqJj507i0qRqBL6RrHkyrDkVf1/TZiw/ZdoVUPe2Yc
IllKk80P0VSl1ZfV7SKzH8kKnuL6LjjY6X7tNy4zljayiThNb7D0EqMihSi0hk0WsPQt3tviYoak
M0WfLnNgrcJn0y7hGobPCduVSh1snRYQUFYBPOqNXmAuZMKnhzAuiwvXPv0elTVowkTB2ec/A1kb
8K8+Ojtpa97s5iPh+Szj5zIA7EEMDulKhVCqQ2MXHqb8CY2HaRRZeffiTByqSuID/4nBWBAmNJeK
GmKvThrfTCer6CiHXs/tziJj+T93CLErcfrCVrLXUJYeXgPKq5CSK5Jkh4qvMqiKtEWx8MWAb13Q
2ZnjWqeW9Lmz7PCQAKhnTTzVevKlXf2okoAyEy6iEylHPVEGn3P7BamdMGJ6QXk2BYmbcEVDUOT9
x/U09O95KP67EetqeKSVHPyKhOWwrXhNf2IocxaAuse9QDYrJKjbEmNgD3UqZDWeAG1WZdONKw58
tsiSN9WPnQeX9b+ymd47RgoM1cCaeT//uhzK16DMCyZfwNon6ZzGgVD4ugipJr4nMUpEivv115PW
tsEeqAlIViVbu9iLsoRsF3EqHUGyjRkYk52t4cRcvklDTymXdajr3BU2hbSLGGPgMauu3OjMZEAe
e+R6tcnwrD4OtwfVtXH7myIK3EPtR9T1JmLaQa75+6lFMLE38+0LAjLtYZLWfYlBzhnKC5cenp2w
NjP+rU1wycZWDXzz6yMlV6icrbTUe1uy0bExWyJy7O7osGkOxURiJJF+8Lgp1hBXsxln4RDwQ/7k
P5fbBIQaVydK29ST/kpOcKy2qHdF4uFxZLi9TCWBBZiMBLwbAYP3aYHaFz+C1dqwNfZYrk9HZj6e
6d4oUVCba5od1O1xutsaKFtaYWqO/wdPwuujkt6+fjpRUM2rajsFESi+JPt6S1fF4vnQyYniIpyC
XXBq8iMgM0GPuVfMUORZ9ZK6Q2mPMyI0KFbF3j+9yr0cYcIDomh5ztHJv93hR0xl1wvL2seT7Pdf
+OVQetRG0OWstgnwiP/IOpU8zHWh/Rlf3yzyTfVCWiWsuyewQP/SPzIG6atP1k/87Vt8oXd4Ty3N
BZzVKOYjC6fJA3st9232CMRIdRsT5OojIO1/oQSdkTD0tlLrXw6wVAekqT2htKBFmv6VtF40jaUD
/xzJ4Ze3doD176WjK61PgsoSR6WCo5fkPSXLTSWKvU6jtPyL71XtzuQViAKyyGzpufPR2puM3Wmq
BhRbhKcm0YaAs7Se6sTDS4tkx6tKzfiL+cW6aKcmL8pdtHmSfIbYbZRiMEw/ZiAGakRluLk1ZaWJ
73MGeMqJZg+TLqaLUqgX51rSnQ/x6eSWkXWr4z6vPUDzJPoCP+wCovEnLiAFXYCK0l4AMGqJpUeU
QrHz5pSrujJgHji0Pa+KgCTGRHmEdm/ZNt9Sw37v74KuNQFBSOJDTxCJYqBMOl9/naQH5r9BJ9cu
G+jcPoseZbLsS0hn7LgkMpQf5Md0wfynSVncph4rF5Xvsnj/7Acj0T1JWQDF3p491YrxA5DsWbYw
U2RGeaF1DP6T/EdqJ50utC4a4SdnkJowci6E2sJN7w5K24DE11wfsYxwSuHnKRdaBXMOq90KnAxF
lWSsGnjoYKmsDuXzIcVWsisCYR8uxl56CLnulY5MidxWu2BlDR9iwCiDbiQZapTT87nf4MsyDrUv
/L2fAXZF4y/Y1UMiNAB5ZPDRV4AQAxsZSa2mRmoeVo46norhpXunw88WK40D3uusCeuPbSfW5Ama
nkoBtDdxwpVkTMp8sfT6l8xmPDsiPUnYNfx4mwPwWiiNL30xRzS04ZJGRK3/ba9j1/YGibpSskQF
mUmki+isLvqMQRYZDN3j7p8JG2lGP0UeO37dTSDTEOZgi8djlqMeSU7tafqlTYwROshVH3cQul5l
cOauR/0/NGFIWWWe7hPi0xVyFmW0iaNn/43J/LUe4Uer2LvK53wE25cMYBLji2vaRzSTM6kS1OIe
wdpIxGuvemxNgNQ0gBwsPYduJ+XNC9qizPU9gn/4uCzGX/Q3CpF4LnTidPYNuqagPvWJ1m+sFpHH
8MXL1ZrjQCFNBWxxioGa8ixf/vOdRuhq0KWg6bm8eeCC+5RSzx6m3SE+d8R6kYcLHj5JHAHHi6wC
tOD0DWrndZI2RO9oi3c8NEQrq6pp6w6O5QzBRMzKbaNqAzzmPgNab+DG1QzIvyi1BQwO6yglNYPA
5Mxg3oK2d4rzAPwmLigKbvlauzqo3AjLRxE25Eagyl4zJxboKQB7rZ9Ss1rATcW54TYD6SlzZzFK
BnPQ1I0o726WbrvpBdkR1Z/uU1VHQLS1xTlUEAdM3plv4cZ9cwRjIsRSPjCzcrVwb6wsA0snXSXx
AjE8jvwGjJSaqpucAwGt/QWAhm00KBMaesb+tAqtPWJ9uJp1K50slWEdTkfaEVLrMif2oflWZEJH
lAj0zAKKQjWoF/JcdGjODH71m7NWZoHYMigfRuJ6kmOsW4R8IpeHLl1YS0ECu7IJCRpbEcCSukGt
GDWhqPIz+zLmarDBLtySFSl+pg/Xx5FMx5kn/k2wG55++HVeXZQ9s6lfRJbnZqNunaKwQNuhUTCE
8QfVnoIBhZK0QutIeKZEqsewxwQeom8lzrOwwd25K4zaU0J/TbqbefyKQ/rhIm6cCBCQmL6qNvyN
XsbgT1vdYQQWyLDoGBOEucQuhbPOX1yqmg8QfMeX1k+NWN83IKLZoj9Jho/XlpLPF1nKWiLsdyEI
E1KLbwairrsD86jleUbAPX32Ixx/B0VmfjwVeyDJGbdusy2AiratyMiriLLHlkLpbL5D6V2uoyGd
KzDKnHUB4VL5wTOZvPWyOKQ9tK1atsq4MB4ZJRMWORxEQQ5Bemc0rIMcXKOGpP+j7bTQETEqFgO9
TvTq7B7M1zwAZ7KToLI++6cp4E8e8/jKNSzZGAmuU4xHLKe9ab0UZ5nPYQMFH5g8zUO02u2DeOdN
pRJuMc/CpDDRkyit1ZYYwb+6xAeZKUMVps6e2GTd4U10lgtzz6LtXJ9vJ3MdCfFMU2bgkS9ba1pi
X5sr4jA/FNb7SvN3U94otPFyw48TiDn/onhXdRT1u8SDkmqxjVbenkxo70IFvrkqxLwpEaU11zJR
JUdEWgwt2vGj9ZqBRR5a8bTE5CwBeJUZkFdPg36Br3Q7nvKPdu/IwSrwbjEx4qo+rn5a544nslsz
gTwCh3rRpfcTOwhmZHW6/iyhm3xD/7rptREBhoCso3Xjnqo9imKzaebncO3MogJWO4Mq+PS/6nYG
kGE14ylKMCMu7qCpu+J7C2UnrzJx8TwW3lfBXYmysGxXvlLlJVY5IXmSauAHTMRpYM5IfbXMXJBI
9CWeKSfWrx9mDS/aN9+K4U68WY3aWdCmP7MQ8czGhhX6KWq6QRzkAO4DLe90j+x2DSpf5en1qvaB
aiSzMdnvV1NCvfcaJBGRoIlUjXnhjpfGQZOdUBcqHfjIbjLhp5xGa9KeDAsAt2Dz4aLgoa5DGOQ3
b0KeJd5LHPFx25W08ZQc9Fl0MtN3xqVvRjfgcNubyGw/VMmAqV7n7J2g/5yCzXs3/c1gmICt8Qjf
onnO6PR5uV+jAaLh4C8VQhPVJ6AjA7kTCtI3CIi+zja299PolWriEz3k9MkERgElsqawrW/TpSsW
bXR66rE7yPLxFWM1diePhdg33C+C5MttmTgECVh+R1+Tqn6iXulnbEhPLcDQpU/4BJuHKgYBy8rj
KPsPWj5dlKE0sxEiXLfRrc0iuZEh6RY8er0c7QnRB9oC9zxda8gMUQoKT0MxfCbrteaDlSyfEn0P
SCKro2duJKahXZB1E+a61+hV99jrP5oPn4a8rJiu3dJor98OAI99rVMGwkKrlR7QY2ciA+VvMt1m
0YnJ2dMQx1LbHsWqOmwud20E3NjHCzNJUN2LLOxXTvEsYOMgVx4SGiW2kKT2w6AQbjAZ3aTuyWWz
KXPwESu0FQI5BsGE8Hv/chxx6Ei8nMImSLc8bfGSs8LgG9BCFP+q9+WJp24fDC2W/Q75LHfdPkcM
E+kI94LpHJRvVHDgJSdPx1aE9lWlilhf9oywI4SeF9YMo+OMxS/F6ZwuUAd+ahJvnz5V/WzeUI/E
owVD0KMaRzL/yquY7UjthRmcxVA5z0B7S9f0A8ahu4+f7KB/nBYnt1s90wYzjzotltO/JzhUJpas
1cayr5hwFdStPRkZ6FpP2j28G74ThyyOhJBkAkfGGFx3WTQIdpKHyTjVQKEE33QY5xBrNW3CEeZm
x7trgVbETplq3935NC1WfJaA5tcavgda6o22mJyISl5ActBduw8Zo+Tyl48WZvIsq7A0K1dM5M5O
ihxNo0S5/D1dj9wOQr1bPsFpBd+/s0UHfBu9IDXDbBbnJ2UCzrzVnB9Yu5rA72RQpaae+6er8BKp
TX0iFst5lr9EI5zJUQ5zeJLADodAOO9V5r3RRFdml6A1POgTqNc7/SLV6pyrothF7FIEqXy15izI
i/YNzAMVmmGB/tJ/uMM5Kjj6Lfk9m+B6gQkm40UqEM7oQcwC8Ze9exbkLmcq7z9g065e8g+YYp7u
nNph/IilvV+yJTgV42FgCzdoCoDInn5K3VaV2SqOyY8lgekdho69UGkBu5JVPsRPt78oS/O+5Gw9
bRdLpngV3Ph4+SbcP9MFe7Qr30ztm3+piRDukOngAWfAD0V4yw0nI92gOFUGnJ4G3+H2ZDKzvmL1
BcsdoYmBb0lvEsQZq5SLESRL9bh0KZDnZnHY+PohvEPcU4f30fVvBZ4Jq10dvRFAqPIDx/9JQFeY
lM6KZeX8Y+vJ3NS0DaY+uSRqlo9oxpeC8IPvbTuCpUqEz8DsUjlR3510Kg8pcIzKPY9DegT29YLU
Yb1lcHNMHYA2zVHIH7fkYvLVk/oVooOHn0fiNpFWySUX8KEXSGsRc+a3fPt9mN4wd9CjXgpkMAbb
Fci4+wnvu8dxNRVynLK27Yt2BwW/RVTxzZA1rlrqk7ua9L2Li5jR/hT75kRGnDRE0uOrksSTU1oV
BfuL+eQ+TVUKiBtUHZisOI5iO7Kq/7UtVEMcNueXK3YP4PgT4Ftm9+EQYNrHhApQzT/2zD1/Gf14
+1oDqbSKfFoC23v872misLdKpJZOQ/B3m7hc+8ktS7jH5nEov30bv9BoYrVBdLbV+oEXWTb/YQ1H
FfXt6jp05KRHNpY/GN1dLslF2rDbLPkNYHs7kqrQ3CIx13rHHFDCAqj9Ssxrz4zp3FWpESBREvWe
rSl1jbdn79yCi1vBQiXv6lU/ZFPpu++XipVmbwvme+ZDcfUHrPXlhHcaoJD6TLCd3mya+eT5EW7q
FOJMTsygZpWizEB/4fh802bHqAZW9vysUQ5UlZ15bdF2cgLTyTiJ3B9VktnpqlunWc2CsOhPZEWj
JxjbB+mtBvm9cFno44zgNZgOhwQR7mvn2UtM3dm4OnEMGqInJrQaRg3Z8GTf36UraQs+ebIRf+Ot
EO2hEMh1ELu1HW5G5D7hEjkeiCiuvlBeDu0Dw+2JzzmSmF7XMAuxgPWAL2IoD11Ms1i0s47FyJFT
q0LaaXABMiumjTcXg2itSA1bKrx7xXND6jjWARKC8KycVQC+QaX0PwofNYILv9KraUkQimtH3HYR
AgAAwYWyAgw7nJQuB1LUijRt/rz9XI+nZZ7XnbDo8n2qQ0wns+U0+k/CSsoRZq4Kyfd3nrnwki90
OeJihEwd68R2tafV7QGlWp//j7VoZnUFBYNEdbM6fzuwSW1RkEbbQZD/0QwMbU3ZPNg6yCuyt0ZN
HVa+hvXApuGoO/VGg229f24bD08L1sNfBZUN6MZ+ELuB1Pv1DsJC0J15PwLz8Dz9CM8F3+x0cHhn
WjlM+lsud64/+ZleLaf3u9tecxeIoIHXZNLWeeweD2TiYHcEPchlBToSY6ZLjApK1m8dr/ynIC7g
VG2/7hYb0J0/ui3ajrQhY8A30LvsaUIUdTQwSelfOg9BOIACxt04gijsNgmoBzTvBxhClAQlpVsd
tTl9gz7/zWho+ZxXoQLgLXJ7UyQpRfDr2q6GuCJlZUe/9tmvUxwCR2ZL9lMgoq/P7s0VozY+Cag5
D2YS4R1dTpiJPQwVoLpWDPPYmxM74s2FGOdCcDdXC2UTIHetNzpK0qyDF+Gze7uBWdfEo/8eJpoz
y5u8aQ1/cFKyZwW7XeDpOITH4kAu52scCAzuNwWF5wQLMjaGbQO1SiuTsLFtnfI0W1M0O1zqTy7Z
tz9R17XPLubR7gsh2V5MPtzR7zuf9KHh/+MoG+UhWsRZjQuH6fh31ooS0TPWqN3gyf3Qmiu2Q+sQ
9mx62w5YWqx20l+peuZhp7MlURgnXxPTHTGvPb/Us8niHedoCYWQzXaPQ5zm7DY+U07JIqGu02hf
spfScYDdFEEWx8C26Iy+Eiwo+hc2ziw7cLnfUM9kjUNICNZQuqFDPosQSQEnI5qaEO1Hyc/MMTXk
B7bZA3H9VnvM17Hpr7dm493JVsJmfj32v32HZgIeRIzCXkGb2Iv7kxPL2yd/cGyGVtFjJu/s+uzh
XQRxiUj/wlDFdxpqKalzAYW5sYycqqKlFRQ9H9n3v5R4edmK9ClEcf+CCiKdQrJyK3/d00PptA3m
n/ZY+sHhetdVP1uMGVwkSjMEYUFVSk8qt4UHZNn3u1mzebQMa5UL/fPMI3FShTF81VJUldZJrzMB
pVUJ0KQnz39fROne1Zd5GUxLAuzk7/e4uq8qTKObM04D0TnGXEWreOpvqM7qwoyURoi0K6scu0/M
nlTMZz3O1MdNEiKBXWxEXgZ2yZt2BwM+mjoAUbxPvmc2P9bWGhRC3Pf/KiCCCL/pfE4hrRchRLj4
2KgJ7MWrC6UGEBNJciO3el3SJwHoR9MuU/CRQ7eDKfvsA12T2VBWBOu7EANIFnJTrxccmJPoAwR1
wCCl3OerWIiHauq5EG13eHh8ghNV2ahykGzMFlDcCWXSpM9R/d/DqtZn/9ja9lprPwvrfVbk0fy7
+u5YDoBu6v5AwSkKXpYiU/iCzfjMP7nBlqStEsHdlUyeH6gC3JvF4+uP4zFDdPFKvNrAo1ma7HVa
Ujy2tGHtaiLFHCC/C7HdNayQQL5oJT4Bwal7QXnA16lVnfiR9IhpcAS2aAGJSBlPe5490LEiGyhY
UCbb47NWzUJcSI4vhrq831e7gm1SBHHsAt1eE8O2FkzYSv5fzKvrNlZViWQiIm8CpEAlTYe8JBnl
WTAWO99viMuyUhk1vfOuLw6h1eq9YcQneEIIwg5vbr8zPzXHJ3nl7J6lmfQhf8GbxwJrfigV3Zfm
TrPnYMHIxinPV+H70HsXCFYsJr34hzHEaAS6S7qYlwWIxn335O5pFE29X+wQlzXERqDrnChBtoDD
qQKnOFHDDo5WsD9pFWq5kKnPnZVEbZKfzVYGeWieLckwLhcSHRpA++PJmz9XXNygc/Yzr4mgZxqK
AKpx0h8VtAcQ6ODSQ1bIZynVhVHcW2RgmKD/FhODVbD2GJ/yMVJiWAb1iC+9ZIykJHq6iO/eL3B2
pOqn3p7nyaKQJseaO6j4EqMJ4yGWA6xBAXs3n4RwN1LNls9dD2I1E75EE87+GkAHMY1tvuoWNYTn
2+Yam2Pe77ofcModSqOaiQpSzPasiCKlD2iY+BkLScq7EIMHGIyKkCmHl4MPHb4P7HaY4OUi7kV3
S5D4vAWbmNkrZTE94ajj4MIer/0mJIszrtGaCtCbMeKYBLcuVuaWl3K1wzC5ItZWbzEBxfJ7bkQk
OF+2Nb8gMsm8Kr9lderteDrm5aS4N1JHcGEMGb7jL8HN+LxZups6GVEWFhCU8+5UwIv7KliYUiNy
3OBvIHE0HPs0hTp7YJDE+GFwGWxdnm7RFTsuDs76iQEPAHSLb1f7o8EmIIm0e3NhIQthybxZxWfX
ox+BYfuvi6R6A8lQz0SFXmhj3QIAGl0DXDrez8z7YV9byP1wnjHRNKjUGso7AkBXOfwjwTWgOeC2
aAi19rg8rvxN5JVJxxdNZAAdfIhA8YccBRTdL+3rf9QUngymCd/CHRQSPjDlwJnoE4cQ2Ymmpgy1
JpCTDi1dRxhrSMZSsgwDGaUlWpVdjYjccK2FHlJqtkxaU3730m1hIMBAH2x7e+7/CYOQrJviVsFD
pUlLEEau3xNiJUshGJVg4X1PubrEgIuD9z/2KkEHkLInGoDTzoZbDmXsIyXds92d48vIWUIqj+eS
DUkp8aJGvHq2j0CPl6znlGycjHBgRVn+Yr56h6eFW+43bAg6oblFp7ZaxtRgmU1HcQWitm67m8hb
0bRG5ZVcs2/5jXf2bvAZT02q8slNW4lrJOpl7B3500zyOjf9TUZODmM+kIG/BHGxnezYdSHP2LKg
Fu/I1XIh0RBCVnT1q8qlze3/vlsPERMeKgQjXnA5OOYwBKt0ib9TH7xkRxLBRNoSxmDdwoDNfP2J
vYiMal81ca0CcEE3E55d82glvnUQY9UrNSlvLY3LMlP0BemTsx0/ZQKl4z6nXBrkrN7ujaStvq7p
Ux+arYf0v5YNSkMNEpMeW4JznMNK6EEn0fsgkv9AZ0cct/7beIJ1VcwQanS/izw2TRB/mZBg/UsI
4yxWTCkju4kjtmO3NUZceacnNUdyVHr9WMpR0wwBwD9wfPD3hWbLrcmRmpCwyGVIWwtp/25Wt0ex
EGCDvIDOiFUjdJEDdLMe3uv/i2LrY5t7U1uBB06logZj9zcSNxLdKh4KktrB2+ZCSKqALiJBp7sx
6S0I8znuUeCIA3OLXLMVGJWL9+c5ulibxQogefFCGd0qMW3/WLllXR8QlTXyvWJ0oG0jV2XOenLP
jeu2E1bf5Lw4VwREG+RRQYftNghE3B5AhBJZC7I/k5+y8pFr2Nhod3OOty2keiDXbko1Cv+IH5xm
Ksqd6dPAg/yCP30KTDoN51CSbX927U223DR33AvO9r2I3QkjjS3M4JdoThSMUpWQclRXqd7q8FOB
TuMdcIrF8L3eTH4DdzVBK0GFL96MBr4vWWZF0cGu+8HmnU251cvDr1T1obsmTPZmMY69zzhbnDfu
HQQWMMr2AI7veRayeVF/v8DvZK4gZtJupgFenEo8jfsKDdgaZjO/biO+lywP8IMOIzXAoBtuaxaC
EThK+jMFkXnEo4lElmA3ldVIk8MmyhCXisu8bFNe+HTr7gSjHtb77Yvgr6DsxbAuvdjHOXj0BcEc
22eREk1tNOdk0ing5F46sT5OuEHQVDnhKjPtKtZcsuU2EWlyiLdoSadWLE326geNxznvZ4FkR9J/
GzH9+FcWXJ9PK6cgHf5UKoaqlTj4GoYxids0r81uhkOcVesOpW73rayhZEAiVgRo2UxX5GcU8VS/
NLmUfuVDuRX/57SCqBi2SZd3acUtN8TO/X6VRATAJM7gtZ/Jd9ELP/IxRZ/lDok1fqTGI1voImxP
E2RtxEgqqjY7MvcJXvRXKvtc0p8TVG2DQcBdZHTm2raYfILFR1cknkBcmLtvPqiZXMCVEWkAoyK5
w+yZQPymQGJEvs5mbSJ5Ce4DSA0t8gvWEEhWArwvAkIaNGRHXiHHAshRx7h+HahYLd5JA4/UN4IA
5duIcKlPGIOgqZvCmNnx73U57h78CQyk75LS+f2BxqZV7NrreqkKPIAUQu0/XCSTS5AefLY/YwHI
z6Cru1RopcxvjkcJbW2jF6rmYT4oEeCRMObzlL8TbJI3mt87lCgkAe81FI9+cT7v3aYefXKFyzQw
Y0Z25JfXZz1L6RH+IjAW1aITUtXnComRXFFWyo7cPu0Ta5RAsg+hm4GoyZQSdWLZxgG3wCgTJRVe
n3hfQTh9dvgnCVezkv4Es7ONgF3NiD+eDnn5Rcx3KGHQF8GdeUL8Ialv/gNirCOKv10DdOjU+t6o
2BpnTdriXxzgxt7SLV5o1sJ6sUM0GE4rtmbiWxCej2n7IhuR9NMjgWdkiSDafqgMz1omoBWKFNkS
dWT+6V+ikon9hJmWMSN8TK4nY319/wMmoLBp/RRwvAdfidoui7DyqHNlmSDHm+oN87mWzq1EVRII
Zq0tkqnd2UCLQmSVnR/AaS2+sbl5IPrJL25FH4SKW1ICgBvV2QEtZnz5XfCC8XZSOGch3QEzYQ8H
zk5WL5oy6M3gVnPdKDvJJrsOcmr+M1QkMwc1kWHtsW4pBmeM3hDl1RldUv7hPS+hP/9lVU9TrCHg
q/qWdNPyFNHHWd6rYtDir7Uz6P38r72dDRLcSNsgpq4Xgg/25uUeCehPKsX/ETAEHJ6RIuieQEJc
606TXlyyS92e3ADMKVSrVWwPIKAEF4MuEvi77SzV/0f/yVre4a2dCXvnaQ0GVa11yEPeAJs1H/Tc
lehe4SNr8G6iaGK2vtgSu0W7AFB1J+DUhfRCdlC8SBgMInXIdfR94qm2fWphqHA2qqSBcYCCzvfH
aaFLg24MpfQoqIQ+33JfUKaWZtPTLWCNGg3eQzp7QoY/p+td5yUXjpo/gH0TnyV8hgHx/Ez8prIP
tDIVXkDbLaRRWG5AgLhudYZ3dxBA6l/axUBAP/SnWSuUZT6iD6/HUcqhA7icNl1EtG77IPm6ajMl
L8IBjNfyg2dD8SRzYVDg8xv32aSOUYeBWDFIHkP/BvcKWLK46xC6g6GXzHMZT4Ym4kdeukJ2DfKx
fTmONABeDp0HzsPfsdYx45aTlUy2zS5j9odnszOPj0Hpyy86Cny+6XzDbkdGWdRxawfpPq507UfL
WLtt4FiSia8DOQMHHiT+Xeatqk8adTZx9XcIc48YD65/qAxZ5tK/s5N21YE3e6uiRiyHVdbvowgV
uQFeRPtlghqcOdI2Sd0vH/aQO56pK6AEegh305meTVf0P5KvH/ofpEhkow8Sc7YYS+FT/zXKstDB
32+ozh9zZB3cZG6kkvkt6jSqcHQWb0KKQn8n25TezDyQxyrvpE5pJBNsF96nCWJCwtlX0f2TYTEX
PHxelbpW1HGEoivpg2b4XqNvBU3QSKIcc4570XW/QUaupn9tIuS07PnVZ86MF4P7p+gFZaG3PfZ+
VRDAwdivf3aM78MwilhERd0eyDW0OzDrjCaPHPT3Kb+6RekxF7nJSlpjNnjSA3p0vGLhXIEsSwVD
MfKCY+tD+rVCScndkNYXDyS4wup42+t6BPSF3Dioqq6RoWwR5w0mh4fyfgs2oBnlVyr4KPezY4+8
myBU8+qAZhRJuPpfSzZLxAAS6xFegOI0uSQl5saARiI/mn9itvAEC4ODjxnTuZrJnHtgYxHjjVWX
rTqfZW4m5aYrbHiIifU5vYGRTkj9Vrgiu+32/hRdq9AN0UdriNBC3GvaF3UUpl/RVaRqBhN1amLs
OIBo1GehLI1jLNj7YPkln2/5xXJXxZLXUDHUGP7bMNKBcczN8UYsY4U17/POO+USDIB2Ura9/ylG
QSPj4oHfuAN+zQuaI7zSDnbgL6xeme2faKKuL6MteNtgl1sLRniQjybe8XYyUK6wnAFvh2l0apUL
kFMfm4GEOKWpLoZKrTFbTuMPUqatBg4SGgo1C8xPggkWkWyQAaYdVIbs5xkQ6VQ+jrEePP/HC9mM
gProO6JYgcoXqZaHYqQpaohQOlAF2emKTMxYZ8KYBG6+dD6JtIGMPypNOT9uc4MlV94EoIOmVCOX
MBscodjEyt+6SxTRFmyJuRtBqrZEGeLc4HOqWqnOIpHcTIbI6QWk+OK6on63UT1U03BUBEktAwSA
5+6vK8qwewYZ+ZMyJpc0/GmJcgeMmIlRd48e+z1xMZ9nQ+KJDXTle83thHbaCXDnDvui2UMBUUDI
bqZ9+Ets23E05GlDH0UWvpwO+x9Oi3fAuoqr1lsmOEtiMChmjvQ2PrJvexSTkuHbzJ7OD1zYDCU/
DuRzl8x9J3aS3nSI8Vdf4XijQaL59WloV6wIHmsdQOPyqzOZzzwdzDhOf+WA0h1w3FvVfGNR8Oos
g14nz/fJrI1OirHVUr1V1ad5XrjGmkK0mYapykHuMr27HgxVzZteX7necyVSHO6dMLOFJV2Pft8D
mLC7T3Hznu74ZtZd4h5+JMrdAKvRWGfdBaMR1K7OGiUgp4eB1ud5s4wwh85QS+4fJwr3NLq4bl9b
LM5feIrqgJP40orOYg6Tr84CpqrH43XwyuXRzhhpsmBEGk19sJbCJmQ10fi49w7BQu3UGY+uUndo
H9hTCp71qbm7A/NiKjsjxZGHurXvhq+kIBOT2EGYKJGWtPuf0v36wko53gPIF7MqXpAiEpEe//1r
n8lYsIzvQMzdbqr40qekeQvAxevzDUF3bBT8vC7G4s4RXLJpZjO/vTMY8a5FTSQfMei00z2+o0dx
72kLQ4BBuT9LQiuG2gXdNBtTaRhs4opu42oRCEBCCW6s7KVzgjN75RQ/Q6PHEVTkj6Je5sb/0nLo
n0PwZhSkSsYcKymVV9L9fWM5VA0IdtL9/gG8FSo2BhEqMxrp61iQMPyfxK4Y71rU0sxJSL6So+Yj
OqLkuYb1KZuIaFl/v8ZUFlpzpGZiEN14XK/urv2urrvx/XnWAmhi4EH/6xe+70YxNLCNALYTDbUW
gKTXTtv7ZnPkV8c2ol8kspJQz9Ez1AfMcDZCc6s9vQwhOiyDoUaTlSO00ME07mLVj4Ub5hQfMMtp
EVBCm1QDJzo/Kkv2EFaJRJ25x84eDNl8pLX45u3c+aCUvv9Jyxsl8fy8JwG6aU3+hQo1Nsw1aPG5
301JgnFWO/UieWraNg93l2KEwF/B5jencaPmrMDaS3PSZZ0YT9Pj8eJZ6fW9xiO71vW3g4dj7Vxy
jDz6hNVCw5/msp1UqSU7jQ07Eut5xaHcaTJESpIPTwUI2nDoUdF/cCil0zx5jBzjLVStjV208qsp
JAacsgtuIVCaV9N9sPbgd5/rF04DTjL7d1Awqhm3WK4zxfZZfHjMJUdH0qmytpdn6jsT8yBO/Wfe
8/MI47Jx0zuNuBH0gi+ZnuZm3csGyJ8f/GTy2mbCUcSbfFCWQNUDxWvjggrEigd9Ia2VZC45/LyV
78QFPK9BhYsYmuGRKsKhMOmTbXLB5Bh7K12oPynwr9n6cU5X8E9n6iY2q7YOeXbIx0P0pUeDEW//
ewhBD3cBfFTMpTYwBKygtNOWPw66JK5MaIu9KDBi3oon4FXkl8RuDRHmiZqEhJeHmS+K+TEgmVyh
aUaFeRv2BxqzIt7eFNVdHjHthYXdVviumFU7mtOqMTxSs9gNO504mUUQh9GVFiUvhDHrB2OYDkYN
aMZ4mUtqJ55pkINFD5FvK8CdgzJYvP+CCkkPvPbpRCqS+VbsbSsjCmj7G85Byw6Hsga35BoBoSjv
BIJ+km6Y7ZOqPT/CuUx17o/WQ0rvR7eSHOBDvgNfpNtuu6TQIja1olHARvDpc4oIUW9KS0bP74q9
1s1X1aFtsmQCjmAyUSAmKWbVguNG0BSRbwVp6sMRYs476Sl20TKfe5IAZ/hNyNQ+4rhJuuwo9onY
mSMI55GbEW8CviouvZa4xXS9tYmOXjSK5NJSvNKzRp+/I5xNawOWmNRWhQj5YAv6FJc+/1wU/xie
AWihF78QBFxzTfNDy04tZhlJSvTUTY5gRY1HK8DiyAt5DBIQERcEHVQVdzsn+oJ8/GnvnN4sYlz4
qfpkPIOgjfNnmMxkTNJz9YcsxJM6u4y50YGLFAOZajDKyx6k10Uc/59Cw7FA3pb8E+HKAHW5RDj/
hs9W5KadAniJF7Oa8XuGaLrHQ1QjwLCj+D4z9cb2Mev73DBeaHuTNutaI1p4G4mMDKUTTU/tsRTN
hllJGSssQUdGig6+8zQjchH9Mmyp+OUsQX24lxSDNJOBbMCLMdigl14i6LLTIhg/yklQdY2kjzsL
PTo9w9ilx6k+BT0uRJ0+6sdeh+myGHdJtkc68A5eR0aduT/muSf0CIJ765D/I45Sbn6fEmQG6W3V
eVfUlE7GFhq3g+dXFGZfrchQUfB0bh4e+XWw9r5vO01wigJvQZ++NxeKiMeUdN6tjb+8cv8ONPWJ
6nsa2pVtBziflQbyF7VDS5PGLKuxq+wGvV0zGS5G23s3e6TkqdaqsstKwK6Xlzl6ztsj56KhZAxv
a3onYrGpS6QV1p9edUoOU8sd1V80e2xTpGm1LIu7ReL0LWrASMtUR+Pes64bypm9kyDLRiHWI/Xo
gRxXNkYwH2t19jU1tCdbya6kYFxM5X40A+ONH+/gAmyebhpKNM5eaT4glitY1B3EjJq70BYvuxof
CJLAooUMfHn6eNsKyVGRIXvh2JB/Vyumg7n1BHRSyV2sX5Wkpgu0F39OYB2xFtRAOQ5x0Ytevn7d
OzJOOgC9dqNejlDsam9E1/b1qIQoK5Z6btaoHUIaR0fo1c4SiEMgD/r2Pcndhvv1G0c/pmK4goMM
1RPkWAFf9z4hVfxzH5z5ckXLNbSmYdvPYHJD9HIrNa8jb8FSTXx0hgDd5UNaY8xn6P7XQySn7Ug7
S+igQAefw9qpBUgNBWfOJOsuY+kmjehjghlUSPx3NiQQwEOEeH23lUDKXWpXSDkIUALoxbcyCgud
NuWOg3VgR4ITuzYJB0ol3+OHrYqM/PHZX6l9E6ZzSOn0IPaRkUP6pzfiMNGme2hX4kE9wHlT8lAr
7KzdJsrcR/ZEmtxF8c5576dtIwPexMB7w9Qm0eOWTdJXn/PaPED46V7ZwkfaybyhfzyRzTo/7NoP
Sebce0DjH9qSCR4KAei34A9yvn1jrHt8hzy0IddJAAY6fcMnLSpX1OFW7FkMek6DZjIrMc1p61z5
hSKBEgefSzv4CgIIKjcAdIoWB7HNcjaasC9a2DvDruPKkhZQXAilcIjIR4epiOZCA15o9np8u9LT
9IcylK1UbblVT7MUlc41mjpktq6INk2yGzQhtW+4hT3p0cJFpYq+duSUAYv1aXpzAiYcQzm2nOuj
RTEekAGJevQk5qaOr7NAg/lRbj+I1PbE3omwnd6kEFjG1i5Xt19BtseAcYMLoXJlJqZwUpqJk90K
HK9hYcLHh4Z2flvv6H2URQ2lcEc18mMuCmRYKeC60BrdohXKYIW89qzfMurjyKGX4yMOfFb+WUGW
6WroG0pfwZ1rmQjgfX4RYKYWU16dBbg5YVfD6LGuMw0vE06JDf01vyfIDxCWhUamMzCG1PiFYUtc
oP/aeXm4J44euhNobtL+fPFrEQq/ef1+LNDiNcvB+cxuM11Sd6JEBmGR7S9ilPghVQB78W26obS8
t18ppahWz7bEFjyNn5FZHWKAXMLcP1k7HZDsf4n27nMVSpIolkR8c8TDxDhyK5sUYy9X0F1MLGFl
X/DUg+wrrh8M39rdwl7FQYvRCv4mhLK5D4PnlD/J/qkhGMXUrI5J1Z+aS3i0g5Piko740STz4FQl
xlDZ34ZpFBTovyEVbINFXc7Qfc0L09pXoii4hf4jPCJ1pvlO5gqp8vvJwrAzpqSabPMLOBNuv49D
t/XgeW4garhaFx/EHIYa67TJiMPeBtImInDg47ti/Qto8nH4RifQgPmQrSrRZRq+Sb0dBuxm3PHP
1OrO0kwTaJAW7YVpDlA689uw57uhNA8uAyblYn3F2LuyIILUWuV8hMAOGiyIox9CK+cs0C090gLt
JJrGepIWSWcm0LOAO6J3WEE8lp7mK8HSvCFJsJWSJxSKNdVSD225cH3b2nksiHWzS/hu+SLCsq0m
ssZz9NUfSLHi4A3pBl3ukG5GZS+7vY8TJuyweiqo1Gg1oRmqcWmSuxhawr5e/TvHCj7b1b67os0+
2AJTP5sYRFJxNcSz5qMNECr2TFr2VsIXzYXeCsbSQlBqro6SlrdAOuy7ggAjSIYaGaC2h0zFNoH5
93WIbcvNCHUC200WnBt29OllMgiH8v6Jl9l9Tv3g8o7HhK2aIXOywz4AsNuTyIyJCE7rtbuf5jni
/n+j4+ULHL+LCthTRR7jZHujom/VzUn9mvSbxdEitp/1fs+MjviZa93xApySNvWjbsTTn7T2jC9l
QCcPBaUhZVca2hVADHebGUZCyIabNs4oV2jsGa/L0PZh3icRIuvxRorXPkMs5XFt9XB9+oCIhnx1
9Ivpgkq4koNvqEKg3LuSWZi1NyQOAW81Hnbxv8h+BPxhJmxkujGe6M4Nh5hmsTIEXCA7NpEQHtCY
aU+zZzJJqxjiQNFK0xisvRi1aKttS5pZdSL291klHlOau3yd1DkY0bn1Ui+i/zkFodWSfWcIvhme
DNkX4gXLA7GLRPyDH1YjMn2jUmgOmFq2U53FCLzBBotSoMYMCCTPif3ahlZV+i0dSk5fAIb7OPMr
0ZxCtY5ekfNVvY8PBYMsVWOlCvwl9seJJnOMpKLm68rmj/gORGP68N2pIbYL8zt3TY+I7AzPKsU/
ulIJHnOLcy9pluUdA4JHv0rv5KnbGq1nbVN1nNZny2zmvSe4/U1eMvfMTAP18kK7dpDTqY/4Y8Ez
W7c3AAoSgK0/av1Hp2ZNPtv/SWIZqhBmpoziOMJ7yECBhYA76u2ywyAADT1/Zua2yUm4uuDWcuaa
HEHFIL5qGg3L0rKlPoihnnE0nWG5Q24J+yY98a7yYP1kRDY/hyRCAd+I2wh6VvqoW1BJYf5i+dxg
O3T9cEMEodayFPf037iAD4ef3PCJuGW8YM1pMI569rQhZo8k9sC1c5sSRtmkkymZm1g16BYCeIOK
9j8w7XcDSgzfRa2nK+Yrb9XFp6gBn0aHStxTiNZroETdMje1w2lbLuWG3A5EC5fgy03d0oi35lUi
6u1mUKM3LTvgL2EEy6oTGoRdO6QTdQ2Plj819AyY3mUDBP/9efdFNifyzggXweoISJCcEvV4iCou
H2bLA32pz6IUEqSYL3eODbRdDX+kIEc7TrxdfZuD4H5xS5rRTQLsKOqnCPC0qmJJtwJLMWfttmwH
Eh/dDdF2OFDt9U8Djjd3afH7uF7BQsL4cKzQmIltLpA3hxK6rGcU9qcW0qjwy0PANos514CKYFrL
5VULhOVssAKwOsOXmG92U5A5lQab/vNGwyPftgn3+bT9SGHILpcebNN4QbTbuGSDcIyg5E5A107g
DOzFZweQwLVfRqa5qDWSz9uIJrc2VPnbJgK5ASqE+CzPibW1Z/zRvplDyCcuRollpBnBf9/T9oV7
+uDtn0u8JTMfN+7WJa3GyDTwCC/9XQniWys4JAa4fgW1Q4qrhe4fE8HHU91fK/UKaAl1r1bLvJV0
/rMWwcuP5FWRuomNheV4l7aMaYdJH/hO9USXtPamkiWmC9JSmSKlkDY0md0+LeUeWj7iN+afg3I2
9g7l1bPUC3lD27hQ75QUy0T6qfM2rniiauAXvRSHw+yBQbHBuAeJazCq3lI2nX2dUxpd/gv7hTbb
qiLTO7eBuPP+ixxt1Oy7tcoaHeFVvITr4VCGuDlhkGWfduovkiXMrJUSqsm9kRoMU2dfRqQcF4Zt
0ZZo1DBQ1Zc/P1U8L8yIDV+PSVfalUTHB1y9IV17XMTjA6nQN/w3eLdLduc/SKhKr9zFEf+0mskz
TGDOoCT6Gw/aURX1qs/uncCIIa/Au7n9zxWeOBaq0SF3eZxlGBJGMB6x5EuR9aFphYA/Ktyorsvy
hVu08ReviYmEB9o/HSPXAVyZZb8tZFAQt/TO3E0APGKor6oNOd2MUVADdvC9srb9J2dEZ62ntIFY
AU+tVSCNNFWPMpcyuGN/kaeO+Hee6v+Jp0j+Aep1HHrCED8qadkUi3L8qMzYvFLD9bxzR1WKRTA4
Rip2m8Ogzeb3xkEKjuDVNS16LVvMkpZD7HBJmVZBkxJ6FMFVkPXAM2glecMPSL6Bx8x9Si2X9Ofd
ZkdJXgauG8X7ssS0et26VMmvf4rFrSGfca224qtnSe5NBTdiIEQu3nWc6XjxtVI1nEzMuINP8LuB
xPFwcH58ocH0UHSXUBzJ8NWnlfVfDCzEqzll38ZWZu0b9BWcBO43ODueO9yAUjlgGMsfqWDVx/cJ
qvMdDUsgo0oKz8J2UZoI+r4mA/qZVzZUzYt1gNpzNczjoKwC4bw+D20t9quJLpPral6HVNtOYkrz
z3ab83xWLebt/jWJOxrRPL6gUM3NRjNZlZFWq7/HAIvtadZOx99/kkg2PCsOvru5RVV6ZavK0u+G
OzS/6bjcEjnK3JYpZUiBJBuLDzy0Yjx89oFc5jj/+jy4wQd+PqBhYYNd8j8GHnVtrMc6x5DsuR4/
YP9aXdbqTFIWlug4Pqs+2/n0U1okMNw9Zay6OgnbLgsjCt6RBxtv2tKu0uPVQT+8nFeRF9nLDhXd
SPGrhG9eyhiZO3g5zieDo2xxkLhUAb5r13eTkjTO6N014xWn2NhQnR20SbcVz2Toja6SGLjsTGiI
x7Y921KBs+Z7wTmRM86oloQ4MG5RGfO6huCm9N8XwwWljaENtu5fqrvZLlAQnFU+1ViCWlYijSjC
xAXZkCM89oQF7Nrd2aoMgGILT4QOakJPBPbDvM7YMO8nfLEolLQ0sc/FT7y9c+gCRpR0HkITnMsB
uLOIkydfRGiT95EHII64nEGNxrXkPdlnBA8y54/TaCSVh4hiX8Mfp+9axqUlozq0tA/JikbaXDWV
+jvNdoz6zT6P64ydII0/lwYR+GL3GHV02PcYZmSCb6eGx33sp5ETqdxUZ8bj1cJ4eEOeM9MYnTon
BYvsh9EqhxDuboyu3bz7C2txwt/OvdZvMAvIhHmbf+Ko8uUtyyFV0JwF5edc3RTGxHUW+z0eDAIZ
VrX/aVvMbgfop7ZsX2vylJ+M/jX8pNlrtKleXwj9bhztikP8ShRq4guO6/QHZfYlUUzeLTVXNDfN
9XtPStGO38uztxXMphItd2PNiZ9+vs0t6yEBQnt5w1G+Lgnj+/HVprktZ+Sa7UWGoUsB7OtkISDM
Sv+U9NoS/rwycvxEuJKhW4q7jWOzhwZxbOPLc9Utzvh3nY2TZuZudaOtQztXj7hr/dm/4KQepRmo
bS8QA3M3k6ib+ENmQEvzgCMicwcNJsaus6bBz60TdwZht4aWlMTC/QK3zVWMvlhsPUHAJa12AwEm
oXpwG8m6gInbVy0R9wZDLax2QzUn9ou1xzK3zXW74xFKPSTnJQl0t/ec7MylZNgxswiPFEjPu6Ht
6Is2gpJ9Ri13gGd226VHN5KLN8ReuLp2QxVW73BVOdyAuTsc3huMtgXjfyS6kxE/oR5WD2q1XUrI
h8LVNqil8Az5DaDM9Eo4lpteDrjQ53TZiQMQNqvvIL0Ms0HT/ZF354lRNWSBUFs5kujwRFRaew8w
1sxFdK9xD/GtvR7v7LYHCtgo1n++8LcUBdNfddtbRk2yrv3VwHbZrrREpgqiABE8kyQx5jTYDJNa
ytZMOd4qNr5YOZKcRyY5Vsh0IAMBtLadcdEf5IEeiFdQmYcEeOpelN5O1Mbo4UrnMDVw8J/fuG1E
eUAz1bJ4T4TIAEQGIaFJK1LW4RyJJ2o9U8bDHFIlQ2iBbLj7yg2oyT7UpRr1Ga6GwHRl7BuzGSfF
V4jLPp+bX2LVJZzI79cPB7gStqMJCzJdAfg58S8fne1NJZto3Uh7azQeZqPT8O4rnA+oHLgyTpns
fx2MNvDNycCypRREyq45K9OyjNGKaN14J8OxcObqiTqkWRykYjm2q7X9ypAHpCU6NUYoTudl522U
TZpFHelyAtEa50IiMHfdSLpo3XAvr8pxSSlbt0LgoKJoDPgXocTh5eejmI1lHci8gng73BJ61KCB
zT4QgUJ6gWuPMxz/Vl4ycCVaya4iX9wXNqb4pAN4VqF7wFRVnZOcydzRzE7mozn61h6m3lmmwHH6
EE9MZ+a/m25Gntnhyl+G0F/eIg6KoMFJpS6QUGD/jpKgcOKMb83d3A+FeU88xtbGCV9HqgTYLzpp
V4FNxrxceAIahPsUMqXLCw0bLS4LQFIiKRi1LwXwmlhHTiEmLn/76BYo5xlRCwWeSxJ51ivuIUY9
AJoRhPtAfW9cMDpk+QAWlRuNZeBJDfy+7didbPzzkhxMJimz4uMCLzwYoZWjtrVMbu/owHNV7bi7
OBeo80rBdMM1y0wYRQlHBLefyit2isaJeSjpRkIoqkZYRubKxxFlFt9uwNvKb++Gw12fQMH5koSC
tOG3/lz9vRByrZaIYhsUWgpexJ7Pphml2nRc50KpDeGByRigHkHcRXIozoo4Wly4MxmlhPOg4mTQ
Zg2rkHv6bKxEY65ZjyL2L5bT6VgXd63Ys5d+oOVMuBVCVLW5LVQUwOL5GQiEQQQ7sHWsXSJUnWby
BLTAPiF6aSXPy6CbLUjSm5nebAOQRnrHOOz0CSfk0cexAiymwNcNa7oq/M9b/C8yFCWM2uDB1mSM
+OAz90eG6dtZ0WJc4/V6zDrVVNtqGzoVNnWMhWYcFmGuhbhoCc9WNPTu1Iwc5Cp40w7pIshso1G/
N1Dm2tzkLrkBt1JC1ulhHir1rJr97aM7eWi3YRz+FLxcZEtiI9bMp3Q5D+HM0/8fjBtfsewOw1dv
F7hSjSuBe2BZycdHOqxAwwrA/Mx7Hf08zIQrLk/s934QtMo3khEi8AS7L4HjCeL+It3bwhuZNaEH
WDGdhJTD9lEGj1mKYWYphBvtaOMVHAQRpFJN49ylwV20BYBsnRz+6Fze2IJr8zlh50nILskn9xR9
qKGEM2O8JwU4S7hxTgNndv3X3Ss3xQVhAOx16nmCFbEYskSP/iro2soELJ9CKZm1hkHlnCJVXfwr
bN08Zt70qLSJYTYkademzqLaHXOflqLvAdHRn5Jf0A7RGYHvWRPI6hXLDsB8mOl83/Vc1rfXYdVM
GnEz2RmzhqtklKdTCr8jCj2bFBxspO9LBtaJTsned0ZjNGC1/e6oNqllyc1xHZGp6TJMRwqAaAd5
BGDe5LqxWLSSfCM2e3IHDBexDBtJxGIIxAyRXf6jWlx8xZX1T5EKHIALtps1rR2z+5n0Kf4ADvyM
L3vDbzQU4Mt29Q8HcbEzvhM8uZOm7MUXt7Q0DJ+w9qAINDJau5wCR1CEedvm6Zv68hwExJ3JDSFQ
DwRTySYdKM5lafr5W9J6Mqodk4kuKnBDgsQg2itSktzufE9Rv+GixKKoVWv3albQFieg4fQHA1od
h7Dg5IAX+s8NGogjG0QPg0enSNLBOLTAlf1AnIioYMPVelg+S76Pw0nb8modpWM4N8XwCzI3DtH7
ps3z5dTxyfW/ZTOckItaqi2iorJACWpJ6gGolnAW/6J44CFB7nN2Vd6TPMue6h++p6WXjq+xg2M9
OmAn1hXHpe+YliuFkWZNh9X+PZudaEdHwwgTAzhnhqVNEV9/uG3cnv3aRX57nl7xfzG0zH9Y6Jlg
M9fkA7X7Q/kFL50t0sXN4G0YQ390At1SliP+HJdQmXNFdZRRMzh2TtzzI28noi0R9iTic7V77iog
A3ec4uTCIvNMB7D39NJWXXZha5QuphlUxNz2YoXG4UgK2UGCNaxYC1kH9EIeP2iDd7oUPGKCKsdj
N2JzAOw6zjIjSbCWcII/cWGxWOgyFjlCX0ihhylqrqjAdx3m8KewinTYHcx8JrvOyctCegbd35i9
DI7y832XchTSnN5SEcBgnwH9ooG0eZUKUSv4beLGC24CM2T13HdJRMlbZpq9/TwwZUqKWvzXPCui
iCS3CmmQIOfzbnSV6aRh+C78alObCbI4alIt8BrYSUZisL/8rUfXTW0KT/4iAWBSatSMB7pwouE/
E2zKN5yamGiyUxzsF/gtQI8HowekuRruZu4I2gFfSe/EwjgbY5wRgNzrdhsrpAoJAyQ2FGFmjQhE
AxGMbMxc277ISy0O8oINYpyXSkPwQ5TOBeum+AA4wob6MGdSOw1lnkzYTVnvZ1v5LiAHMfR41c9M
Bzp7oUbpVszQI4B3IDb1hAI6s+MrQwcknYFlMsXJXoTTA4O6dxkE/EDemMh9DiK5fmykydlBXBKM
U1zuCuHCwDKPQRoR/nYSftbxS5TMa65feyMNZzwxDhPQGQ588FQNa3ZkYGuCgueOJxDF/KODYmqa
3kJ1KN7fniVQ8tnQ0oGEnjzhXps4oqZMM6iGWKnCynd9S/+O8dYZvhTMhbClKvHrqROapAzUXv4o
/D8SciCaVggrzxZTg5KIDSM/PATdZ8BBBKJPM/K3IksU6xV1r36yzp6wGeQ6YplEh8IT2bxhEwYZ
9BaCRKrfx037jLWuLd8fRUIHCWTII3Yzr9wlMpftceo75bgVxu89On75X3UMN7Cb0G6fU/jJo6y/
8189wDg9g1ug/t49HKVqKOMQIrNJOnMB5oxcyUPm3lsdst0AUcXKY19w2WDqkipmN0SyuLgCY3Rl
EudJdBmkR9tn6zpfkoeBPHzidG1X9FqtSNuhBitSxyepbNpZY5POEiDscoR1iPor2xk2ArwcD4n7
1mxwhaEGafjIx6txfEPBR1GU/xFmMowfqs3eQMSRKJl9xa9k6AfIaTSH4UR6pJcG07Hyd6a3mfpt
RBynFYZcqBy0tAC+gNq0tZtaaR43OV2ZvDk3u1XfDs7EHISah7bVgyX47boqQUCxUAoom6R6rRcB
MKagKjWoJpv7F7Z+xy9an97eOouCimmQBtsbpHG9sF5PZFsDyhQ1x6HzmN7hlTGZ4gESaGJYYpN9
My/o2+NxSUut5hP6DBe6w+TsGhkOUNfTz7Bpwj2pzKJMEISJHxSzUgkfuAUOhfnlaIFX8DISLXrx
BdfvZuuN+TDgEoBV1QRJzaOVVzNpVT4lqQD0YQMdp7iP0aVLfaiRLHmCGnlAyy2l6LuI14M0FiPl
THeqnssCYru5zXJs2TM6bFcEPSHWX+se7wkTmW3BkiGOFWgaY3EZBR5TDvg6mOjy0xmuDsHONTPe
bq35nyNvMsjtaJTFjHgYfceuKPIrTtryLxWjPz5f9i5oWNshdrW68jZJdVMMx1B8Dvdw/fuoltx8
DzsQQ4pdh9t2IqFdw1xu7hwpYsLQ/YgJEYV3W0k2uDnILjabe2m3qAxilG9TGnnKb4VzlQjH+Pk1
N+5E0UdHdvcOMwyIKt5LNYxy/M2pbmCmKyXuh0/XT4owxPEapEwCLX8HSy6DqIFXBVJgRnvRQCM2
FW/0mPJ3zvtT3N+c3QuR8lDPJWoSVVLTgzsfs7oEcrkshj9qY0Xx48C9smP9wX2Ug+n0+7gQyVnd
31KXvQZM4v95Hqin7ysxinQ9AuVfzmsnj/1DaSCGhFuH735XWGT7wiKDVcDcwR5+R68YeKSVyq9C
RRdkvbPusCKxpqEwlYrK+wOZohg00Jz4zEGtxPSR7ClDnJg27lZHij7Q9ldHCcV8XzDtiAEspmiI
3hLz0W6TXy+2pWiyPsXX23wlhyKC8T0noia/ByAv0c/VSeDfDwb2piy+gQNyXr4jK94iAuYabDB8
U44k8HXt42kwPS+Rlw5VxPgiRa3iczfDGB5Bc8tCuVu6bUXbUvBaN42FNqpRgeJQsJvfZFz7mbyV
o5N+X6kC6cVf3Ozdx1fDFaayyveHe+FEFZGwWqUY9Sh1b9b6MdhlTZ+Ed/jVieCn+GYHAUj8Kay/
X1lbgiNtGmutUkVGTyWyk8rRQLWlH+2GiYfcMqtsGiKjCysMzTpw8+q2qNUiudEIfyuxp+DUG30a
LU1oemFKFug8T5lTn/YvXz4mJR7UMykBQcMXEpawvDdGk6YmGgyHJ01woM9WKt7XuI98brLr9tqs
NMRUYYsYZGcPGXN3h66FSWihCULT7U+CWUoVcXCts5US+bSshlTA39h73/PGzd6Wpzohb2QYO/M+
e103Ko8vMA53t9y2Yk4UYJw1cSy4wXLz6r3pW3aFqdUUEszZGb02mpwiXfDz+8HuuZDD1y0yKByk
+MmtPihX99AuuIu7FN+RTakxHO77dT6+Um9JCpveW/tZ6ool0ObNy/AMw1txZCKsvJtACFmTBndV
JIS+cGSFL9gTUiOsEB77SmKbNUzj4uL64FusGZi7xuv/QsK/1hcYiCDrp6diUf73fFxcZKk935zQ
D18rwOnKOrxSw7om2bkfG3HVE/fqgkkDk8QNhcthXhmInjjSEhUuIbIUgrGPKhsDQ9N4NtRs9LD5
6+NvBVX283DZ6SK7YoYok+ljtOyKui5Zg/hiO7oy9KH3GbAcDaLecoHMsL36vnpqmd0E9D7Nfijh
4MEXuOMztlad/7wggplQuKmRWAlhLdLGWYEVDyVAWCxU7MiDFLeAsjtHSWYcvwFE7X/dd3iyHIyt
BZwXlK319RPNH6hIeZUXRktAA14sjFyqWQVGZfITOv3JuDS1l5YIj8qsEt+M0ErSOw95br46yoOV
riT+CkLJIgKlufeHRUW9NFOPKrK78TtSv1nKv7LEl3pvPs41YLHF3UeQd6L8/OhndJlCJTuPttpN
tzp9NKi0pOVvKSn9oQussyG5OuEkXNhkrfU1sDigcng4XGUhz8VVGilnNhbSgFmFeLvFJ1lCuVgY
uaD4Y4zIv1hx7UZIOVrXyuhSQkU2awLq2jcRM+d/Bz1rvSqkELWb3kYSg6vMbHix7R2+aZ0IcjcY
SQEv/5RimclTm+KaK5WheAhGud4sEE0VU6X+VodlMUbD2HbaPk4IfewkWOWO4/J2Eq0B0EHlzIHL
TzlSD1vK5V9kFA419mMyG7qHuopfQehwr5bw036uSs0e3wXfLgoA/djwyD+nqpvabWL1JUjXEPyV
KhnM6kq+4fPmOi1d3R1W6OX10/hzNe+lBXHEQtDok3YKk050r0UjP4mMM9KI0cIueIgYHTFpF/kH
g5HiMLRm0dasxbCynUtJCQmNR+2iwwbNERNKhUwdptAigcOl4tCrdT3tlDYGXMukGGahL1tEK04x
qQk7QVzVZcu8NcVhfxzM5nLnFKPXkPb0x+BPUY0gt1PPmgZ36aLnTz5cXLsLOARId/ZaSh3UW0+g
dp3pz4m+zMfODyo6RrKWP7XCUPpp96ACjjIuGCJMlhaEiLx7hrHNXN77BKRdkgL9r2kGWFmem+au
sph/N+/oBgUW+yk9fNs/MxkREID4XwB9BONU6GKG1zPVV2Kt0wK/1GJ3wO5EccXFPCpdlgGIRd07
d19cNU6X86nAa7Pf5MTGM6DD4c0eCkbxRGXjRWtKARWL9Y4UN97ml7urygG/bAUDULnhdPnDClrP
dxJA+INBIeycmfeeBmoszgZONXrrp+8W4NvNS7rMnaMtq9OqBfTnng6HhMKTkJcycTDVZF6Dqy83
zonHCrQFCa6aVyyzjvN85iGgpz83R6FdIMzNT8mN4CYzuMFWlgidl4zva8bnu6EyKXuZQ6BzHOsV
HfoGk9rNyeW7Pb/jueDZ8g2V1ZzR6e1BT+iILmbjSy0ktGFohsxrOCc9DCu4gJ7sHmcAZgotooG5
WLpMOSvjpMnGTbpmFaqOrx4iECDHtJToj4ni8kTytUW/qt2kMIwd67Z7epVt4fGOnip8qvjompAh
4dQbB3yEgvT4c/kIuZK3k9nzbUuuB2N8rsyv9e7ikBNooNN4zepWob0YSRqzvCMKArtPwZvNiHVN
JExgLR7xd/ni13mNFNt1XVH7CvZFD4y9UeSG9pUPgfFynPb9kKuuNYmToSyr3jwbf5mBvNg5bqQa
jjjE9i8FSCBVGEXuvtmXebnohVkYvGhxzTbEIe4JSHuE7zAgPP+8Q8n65Keo5BNITJFoSyDVOuGP
T6sD+9rvkaIx6Uk0iNBk/WwtYt/KKV30IUUKEKLjo3Eo6g1CxNnTJa+Za+nD8+DEEuqsGYE2JuWs
ygQBN3ZW+Rvr2NdNy+sNg1aYi9k3gI3GeMeIRNmPNcQw0WkcsgL9f1xQULB4sL0S11QBeLpEFuJL
NC9TCoIp5A8PGbQK1gE2JP2iOnAYwtXA6QUVbqLicwA0sUZ0RJ3npAk29FmZu7L0SskuO8kV8aYP
x5baMU4Kvm6Ofieu5Fq/SNuYYXAjV5BQOtmvwitZ8rAeZz++6pcAmncSE3sKhw9ICjx+GqaO7iw9
Vo6ESzEqWrx6gX/nrzZgWT4ZY2QFA19Ih/ERP5bBOmlDlpDMFAA5+uZjNwfWEU6AwUkM8pXQ26iP
v2Avn3vufJ38DmhYXj3M+pto57P7RBuvTcZk+r3Ebz8tEyJVw62mQRjfwPg1B+nwtutKZiIWGgG/
DbaPdFnniEK5BFIX2arcta08hka63yLnzXMBjJd0ul3Wb9TQpQH0FiM2yIHtrNTkXHMsVckCC9t4
qXcV1+W0hoWc31Ky3ra1NXZQosOeucOeh8hSJumxh+arl8mL1btZ3YZJ+ENgFGB9rkNNbGULnjcf
ba89B8Ot6tNXXiX88wzBrAvYv84hBOuBYrTsm41XXhlg04xIjTTVGSd8oPW+xMY9nS5LBieg3Tsv
av1NzRh9VYugvmXJ9iP5jnHj1WMvm8qEKx2YXcCxL10xgbJcVJ8yRg19rjajR5Sscbt2z8BLHqq+
H0u4K+FmZ3Ksnq9kpwD5AEnKZqCrhcJTEsr3dSc56OPZiQiDTn1sLmYZyrViwQiqJJbD926xyR0d
C7J+SpgGwIefPZvuvRRdHVWaj9gDPgMbaucT7EFbgReM3PGBWcu9nnhc1rw5Hqi8AlkMQzX7ZFnB
wBaWgRY6LXPwCKWcdeQFDz5Eq/rKnTpAReobqPE0bSAdq0/xGXZRtS3PSZbeQ+5F1YX3BLwP5Jc1
VYm4KcBgTaz83RZ5ESrx9GWv+76yCbYZDNjKWAQKYEoUgwhAUuI3y/fe2mqF0HKD5Lpd4mHPlxB1
4l7BoVPaf9y1ybg+Ef6D1TP5UMshdCqOjxVwjQJu29g/IUfPweRy92RRnZ1+u9F+/S1FRMHlst94
bVfJ+YTIgYQO9z/LyPi5Bsc6QVoWMacw4ZvoU40mIhuzIzZv3qjmy6xbBhlfg3B3ttRzU7xqDPSr
4qA5jIFvIWRb2oP0KdA3pPX6yxdTf6LWjzpNyBHadOnpu/UUbFSXaz6YbG+wJNplO4N0at7stLYb
B7ruAozZRJhL/uRAtghdFnJBra+1371waTvj+I7gxXa+YX8fYhK6YZmIonvOPyY7ry/AIcRD1Bqy
E8t7xRS/hwRxhIqlxP7ePOGgzhxTPNkvEaWNoxxL5Mp4Q2w8UBKRkQrPZjKCHMhunb/oLTwrO2PJ
fzUU6Hz/TYLLHCVTe6do4JJxGsz6Pr5/CXISyONdX+YIrpt6grLFN/K5MoZpFH2XdXlmKyNE63yQ
mp/in2Avykrc5va4LBtOzHAtZo1SqoYvB+JTEmmgfdDgoz1fK7vB+EpN9a/PAx9ojDvc37ll+hD/
KiVHf8cdvnuqoNzhdiWmiHQmbWS1Er8smLNTXaIOVc6fuTMcozl0Q2GyGEaH6R6NnM5Z/3YQZFNB
Np2vB93Jc0dG6p2LLl5S9oOOZ+yfIBO9h173sMVYJPAULu+Gy2swz6Gxn9sGIp18iKNOZ9lZvzPS
r+jMq/cK3lHvK6GNqZ3IHabb8xvQ5y0mznZ9X7sK47RJcSSSOLkPO3w1PabkDpPi7WNnrNA8XeLP
ndu2Q6B7rXOKKMI4Cp3it26wfDQzCfTwBi3wadnVh4z0hp32396QN9GjZ27CTQqyw2Jc+GZYnL+f
LePBflcd1P9IQZHlDKJuvKrrb5MRIBkDinHZhnTMT3T5mHYk2SE8zf2umvHY++PkVmHzal8mgCsu
YExQAK7lawoSdPJEo8Unad0KpQKxLe/r1g7777df7VokLB57UBaziENdM+vFm5Sqcv+9m2ey8bWE
1ptz0257XTk4UCo/SV3rnMcwv2g/MtW9x6dH4XzZV+/RB8uAa5gpT1jNZSCJM7fb/YRZRGkliDGc
LQ3yQ2seKmXbePw1ILxoIReAiFlu7wsfqY5J3X1bpU55hmdGne5ec8Skt2enldalmp2xZnD/gCzX
75RzvOgXNenB0Eo97e1OGDVTQovUHyIL4E6ZXAOi/a9esNA4zczq7DJk232ySGAtqLnTnWKyRGug
wQ5fRbkDderCPJvyXJP8NUzYoymjNNm7T+SocCafqbBxGqMenSkHdmdoRVCqYyK2f///JTK79Zk7
FrTxQUWuwdk7eem6jmDpHTT9i4SNjMQzJTjvALHyxoWf4pIAyEONY/CkX6JtOKLBaMEWDP1l3nFp
7DXl0bYKngrVpjFAR+Y1PX+DJk11Km4CHhEUHUnUl8V0EqZCYaN3pCUCh+zEvXh2chEl2ph0YawL
AE62nBlAVhftRrybTAEVdVW83hCsgCVPmfgpZXYFcKMzuozcvAMPsQeV8whmDW0Wpc9nXMrtAP2j
qPTXETmspG3ZK1QnKJFIpVBL11ebZrdcoPLaQSxHPDjLpHKhhBt18Cu9btTuMg/nkXW+YauC3Ksw
I7IJfHccP3mpAtAjSq8XCS79rdtnDcFpkflG9+hdZJ1N7d/8lhXM0i4oWWAxDNJT+Q88Lv/5784B
vQu3U93IFfUT/1QdGHRvZidpl11lMT16zBDd6ftHGkgEhN7xgJ/qpuo/3g3ij0j9fMX6FEqI1AUx
rBAj3u8hfVuiWezE7UmZV0sizraxUDmsU6lUznP/pfqWAUviG6mR191jQKDDTfWjlSAxC38SsJD1
T/+kpYMYUZ7dcGtN2EhrcdPTX9LT0J5m/wU/43PNdxGsKyLciXziTFp6oOAecbKopYYchEAPKUoQ
z942dQYqjy9ThviuskkxoMYNDpivcuS5UlGH+QlCpLB+hCYuXV+3XmX4pJWrBnnnidLTyBzOElOG
XI3hQ7EgQjKC5UQubeKhBb7ELGyVYIHTunsqbwR9tspvLE3i8ZgroiwoSkdHSOW/FrAqUJkZVtdP
6a9yy6oNmpYFtrvx4++vQE2E+IkRQI7X4dj3J9+vo7A1WKdACr+ccH8z01QBFJD+9CwIMZrHBKce
bIhmWR8HrJX0upZ3YqkAfmL1VshRVRrTbnUavVKrYPXSAUv07e+PtKB8APucQf615MGajSeXXRR9
VqBWKQgJ3P0xqe3og19BpOG/drUi6hO0XhW6DJzSAgLMcZSCvxi6/gC4sG7Fx/7Sin1AZNCZwhnr
AV6cqfvO0225LtfTYy+FxYvhTYgg39ERHg1jvCLiJOzpYtYKzR1pQ0GuiLyBORAqjO8WXS37R6xm
jAYhWUnwFxYDPGSg6KaXrCgmPJX581Q5GquffxxcaHfFYsMagkB8wTFp+NIrzJ1XUZkeotQbYPgy
FFutgmzsS9Vvk3sVfAsDetj8Qo6Er5rpRqHfUJ++uNmKxxVvUZOO/d04dz6etT/HGRsOlP5weGCk
gdUpQTvh10CjQ/ySsXP8hoH82RWhqgVckm+4r3EoFDNoQA2HMFWypsryDQ7NtYGKhugeTrcyWTqY
g88UIlWxL2Qr8zH3iggD5Nc3R89VQcIlduGJyyFQA+wSmJtp4ZK3VRyyUpOiVMz2Ws6nLoJDBt63
q9xgaFf5/xaxnQaXQXdGkvkcbDY1OoZUoO5dz0HyFQ5dh9418rl/0b7+fv+ubMbV2DA27vo1f9d8
rUSYykWjePjYbJ9uNzhFmrJ2bBgn4jShGKlKmS+xqZIYFKyVgHYqkBPIHdCfqfG9HCyPUeFYlO+c
SUUIkDdH0PTaRZ27ciY8N/DxPGGIVyEQs6pJNZ/nIS+sNQG9ZMsGBjIJ4Gsrgbngytfb4rdBucty
DsEvFfyaAqHFAutmkQ3JEWiX0OxG6T9NlydTi2183hrwzRhF84KV1kCUkNk3FdZtRxF/0BYlFWCe
Y3a/33W17OJzHh24V2zaCu/hhp+8KNQiHiwVGM+M5rxTuuCEl3p9aQTaJjfS9tu4la+bIH1jywHA
xGs8xK5VYeezdEdB1oouFMm8+BqZBBWiZJhdbD0WM8UUuCRO8EZZXqyxoN0Ne0vC22hW4wVnKWa1
VNcEzrGKeLgWDujmEFL42QnJorplF2hpL7mHtJLLsNJRvnOV4Tz9jZQJHFRMKOEOQoympX3f+nQf
IQ6pGTyl/STsFewSbgA6Z/mAYRG96519bce16VfYEziwfQwFeqNwAD0g9vkHB6VEe4naQQQTGEOy
V/AO6I2ujb7vq+WrS7utLXOY+UliVBXPpWhEg4U7BrQjbyicZ5uJ3I3LI6grwmkDb+g13t33grRR
0ruakYx90P21J6Ccaxs65b1tCSSNBafga1KHkaW7vtIubFCe/AVzxvA8mQvrbH5YZt8tSLyne4A6
pp68hPGqDaM5wZX2JNvLf5JIfyi/CEtvzHIpEGJEcNsx9oSkhsPVlXZYtIJ9hWCIkF8yjQ3hbnyU
jDZfPjel4GtuymA8J864OxDjQANTO7N+/c3TrzyMWTH3d8y6+yGTKewrrQoC5ARnjZeR181245Qq
7WJidTBWpR5NNfPcJmI8ayN3hRadR0W0KOADe/35MJ/kAhgW38Tsr6dQ2tHyjVHv3nncsW62S29a
bgRvI1h1UH+ut90iEPbDkCKRHoAAbM7cSmOH+MR3UfMX/CFShZU4DmeiO1p0e8ECmAJKMlLRI7Mo
8BWtpKWjf+RS5TVN5Vi44UlB39lZL/f4KIqrFrzxdkLF2CAily8CRqi9Upw2wisAXeV/XlQJD3o2
4jrVWtzBuqFdbR2qexhAFBq4dHvdR279klo/QquvxUdHB4jc0RXDN70ebUHqGB7D9vIgg29lK8Fl
fhBHxztoNwqfr96IoIwKY9Z1RoCCOrjFbr4q3reF/H/lQqJQ6GRpX6YWs6ZIPnqeAfHeq9hPwkaD
DR11n6IZf5R8lPobV9gVeNwCeXAT8nay8qufVotdYGunXe7gJVldn8mcCaf8nvAQExAx/OotQmJE
DaoVWlyW/cupOVi5307GvkYPB15kNI67LP7GGH0D5lWf1zjQBtB/k/PoaBm7DM3aYyUdA6tbDGSZ
fVs/yjfOMHfztT9afzIX0942Sb3Dr94xnwUdeqBMeva1+88kzdRqP/1qKDeXTtT0xb1UOc5T8J0m
/kFgcrPapO5XaK23j//SjZb9OhRbGcJ0TNbb3DSdKuIwhrk5/BuL7u+4wfEFVnWgsd7XgL4okwaT
3RMj3gQDM/RMyYsr0NzGbt26WrmTjEh3hIqUopdbAutDjzcPTYYQTJiYlLnrCf6W9Fdbqk4aa9mL
gFvgtpEXFCnpYhNQOGPpku9sxppoBYR+rlVOFgpXOY73SIb1fXGCJjV7YGumbqwaBiiUktOb1TgT
H5GeLwGaJ8gJemS0CFhRNhZvHV5Fudt4U5HArUS8mrc7C5Mad9DPpfB/rM/BkEiRNDl/0kX2/6AY
h6a4g9+vO96oh7AitSKSMotRABtN5AqhkyLrtf7bMaYc1OlYBzZu+vHqD5K5rvwQFvhEtOmrCrvV
J/zZQYjH1uLvR3l1SsllBltgHtqy+0fK/HiXdaFsQ8gW9xU6VWLrVyFYc9XahwmU4nGuIhalpuYW
yD1lsv1rLHKy0oFR7NzV/D1qmwqR2YfCR/n68E78rDA7Wp93gcgMxcoxa64TqDBG+0vcy+5D5d2y
VuenTR9EzUiyipa7hsWzw2Taesqb3tvg5gipTEVyXmor6iglpMKlwfSoxi5sV1jNpCzjHutWox39
zlADxb2n3cRrtg62AHQ4X4eC73Gp2bqAYxQZgFkXpWyKQd7d3Wv9dyXg2nYNc3FIk0lTQIpHvsFh
Vt0+wgzkjS7sWbVzTWPS2aEeZS/5tWQm2WMs1EMWlp1kjE6N8/GZ83vsaekbdupqeAjihjOEg6J/
kuVczzBMladLlm5qFF8xfGyRITYsYc0omjs2dUcUuMruyx5p72MbEXPj+BLye+cqUWZfLEQ1BAkb
Z0dp4xqv4/d/SnUhI0wyQglu53nV2Q0SUfnuh4p894no7+2FMOL6egtmiGIdaxDKwvF9WwzsOUDF
Fxh4cGKTU+h9XWWvquA8hQpuhj7W9fEX177+g349G2Wc0XxcwfwKhaeRKuklv5x/kJjajIZqClt5
Fu7sFGSACxW2obe1LxzFGnGqdaB5rSUuADsfATnbm82UWDINc9thxltNz0Yalr9w1tHoXM+KLF/+
pkz6/hKhHAdFgR5bs33kQzRQ/w4vJcKcW7ZPix35bO80uFw7jmf/mzY+9N8AbP5LA6N9ZgbQHDUr
SxepJF/KFwD9kPpthnELnBq7xNm25pC9+EsAFA0fRc/6lCn1ACpfmSAJt6LbpFBDNjRkkE9BganN
YcAhocOxoKcWW155n1MvLTsOipdpgn6qxPVyP0mYXMzuizTCQ3IQqdXgHHu7DkfEhaQYjfDX9s2F
wxzYuKwKyBGlbbceiUMLsZ4TRilwcClT2xhoggGK850SaDZirIfjNdo7GntNSK7M5nUW0SHFY3Ke
rzUZuI1vXGlLJT6mGTcCRRtvarnZBnBSOHGBJFVggx2vgxhMkzN2mtxkFQ8XSCeXGI4Bz1MGyMzX
GvRDgJzjWlZpB1XltyDHdNVVNdvv0OMariVAxHT6IVTmQYHCxBbsg21Gorchrh0cPQyNpjo02x9b
d+qIzFWv4WFD2w/ZLxu1cPoORSJSWxQOpXztTekDrsyzAivMd1Qfmk8StPBmJl5p/dimETxKCeEv
ryCTIMmF8Mk4+YlOnkQuFRhu6s4Jyob4ul9pYeDJsep7uM0nOK1d5LKwUrzpmaC9bCdmiW3jU9YC
q6dbZmFAnCgxO+En74TqoCcTMFYzMWwJEAUqk/JWjFVROg6ybiX5fdDrk9/z+IntdNwWT/3pIBx4
rt7oZvOYOWlNTgYRegtGyX4EdGrh+I4s6ueU1UJbAdeYWSbiepHzk8kpR22JOgIfJKD4ZFQ0Ten8
KWZXN4O9wO83lOugHRB4T4wVt8CaesGW6vY3ip9HvHOtFFpCnSi2poxA7QXdNvnYB+kPNk6VN0qv
EvMPpzCUvZJpRKmLPSc+eCFz2K1wV8yYQkOrAb/+KFNXaV/JzuOa9kFvJen/eIGvwTkkZTMsuh5b
xYkZuFJ8cH0GBHBQkggDBrZjw+EZgxFZ+OKgk1lrUg6nId4OUv55OV0lTICbMZPFqbSWt3/Pumqn
d/PnF1I4DBZoKrW5qWEzNQeEc2SIIFr6lf4+PbF/rYmDaCIZGO7O+MzeEGpTvfClHLBZOmzpFv40
YSGO8DRez/etkaJ3oGDoUy70q86VoH4gSZzVWsmUGW4/PHIoIpVVgh+bR/z9UxBhMlFfgw9qnHao
6oTXKHX2hKlori3Oi+Z4swSlTCKivN6vYPyF8zb59UnMFT/26zSzmRArjWIxJ3rIwPq0pLnWaYmo
02tcUPlXlR2u7dTA+69Xm3ZlcfOM8YHPsndp8N3dkqcuioaCcNMP4IKih3xSslMl398D+J7Vp6Vc
KbMskA0xbYx/E/majtLy7Cp9D0IIIgwFLDzO9RsU0DclJOp3KvsQJzkHVWpq6RDvdix0jE46OaRf
2wNem9YtBKYJVCxjt96Ea4TTUkEPT6LlYdvnYcugVPWmPSu8ymY717VfZ+ykilw51BlsmxsfS2uf
ynokJv/9hGl783CYNFFnaNBV1Y63FUDn9LCD/5olbu43dhxrlYufnWhivrvIE+5y97nRKLcfdeJP
ODGTIXCNSXv/lHOCC3dhqunPUW87H7SZtiVE0XOHhUgR2OVBmGy0X6JTO7FSB5LTfFPWNiuyP3t5
Lde13xXNfhDRw9O6Yh3SupRMU/YVbsioFJAbc7zyWKfGzhYcHt3jnDl5yS1viKw+/E0jPTfRTz2f
3TRgLHYSQ/3QRPKgED7ClEw8ESPanTcJavHKx/VEcDuIXlN7KSKT6sLd19GvitVTt26ZEvC4kIWn
2Gy6P6dR0bkeVJGSP5aFjOY7e2Y8TxVOW93N0LFbzdW5OpOBAKHH4+Zagap/UnNC0oiaImVwhd+9
CFtFnS7crFfRbh8uf1B3MTNGENA23Yl/y0zxtBgoZOlLHHHB/lUnKQVsEWzkCQxpA+JALw179tZI
1qgIolplqPJaqgAer0sv8/cgfLkZNyd+T9HmQ9FzwHwE00Rb2gzsXmKtZM2QVHk22uYUZ0OXF2yb
T5nqqYYadsHMctXbJKVx5mD/2Z9DC3ztQd/VpDHC/yT52Ut+aEyJd/QtRxu4IaX/IkAvMPnpwdEU
nYTOfmnDqzla2VcwijSkgTRh4jpWWiat5rRgHdpSoB4ZswqYKOt1etvwop+03ZT4KErSa3+HGZ3l
19J0izcEbnr/oa84meUqyIybylM6rEKJz5Z3WZyHhoqexx/3176PDsFXeh/PP74pYQbimxoFqkk3
5CBRejvDbthEmkl7DZyiC0GNvLkihBnRLr9PVXOCXup2J6quE5ajfVcnawgXMrwZxZD/5QF6d/np
Iz1cqlYiNrN/uzWOvbLq30JCOiKkXNosgHgj8n5j1hL7Qp76RjZJRf/g7gc8Stu/ojQyD1Ml+Z7c
C+P63RujToCtapFNXjz41f2WthIkgn7+7GDHh3PSaM9LNgRl+lk9YfwprfHMOE50gqmIOe0ZqkWi
oTPiumnszxlaKCHCd8736uO14IAFqGvIWGjiP/euAASByF1nB5FvBvTMQguZfYZsOppl7vfjeNEd
62CJzgev9jrs82qaU8Jv36lVfrIoEJRXmDwt0vNfDxv+2gjl5xJSzYNJiKKbgMskaWUvPQSj9bmP
EgYV/5fdl2P97titw6b/6b84ymnfNcKwqGfoAUMfMCVdojzyC0kUyPSNmX6itiFmktPGq0sYCHfG
xfmzTAIZR9FX5TsuOJn23iF/v65qABRk7snEfmt4+/0103e1LwhvwIko2kQ5XFcDGhY3VZ1WhtR+
3D2dQa3h7niSEFBkrKdTrpYZJcsJvmgngUSWJQJ3vd9Jins0LCqDFfe8TecBqhgR3PmarE8gJbky
kOrQBFJykLZAtgaFCOC/zEXimBJs0qF6rAHlMigX5hERK4Qhr9VAoFgQivjV881Vk20VsiPyJC5S
EfGKWdzSdKFaoQITBug5E75vE/CNLbu0FQXkFMYSohrTKAIT7Y5NJujwS6Hg6pIxfIGk37UscgdR
+kAN+QXOgmxe8qS4hbmpsr+VenSucTYtBfOzAR4hFgx8fIQQKBp20+soiZod+KJN7owsvB0H1GzS
79d/l1sWTp5aZppiIfTpCH8c/AzlDVHAt2G8XZORC2whVG9rVQpsDf117jNJVqJZb9/qoOmsZR8P
aYTTAboqMou0WeLcNv7LFublSi6fPC05+VcWbsM34tkqdUE0jAmZpjbTnnMn13dUbXtgIiybN0Se
9BDq0jYyfcYDROMP7WMa4ydHQAxi5GEsxEopCJbJ8xLyoyN5Ez/x8W2qEgGXqsn5qll5z65WwPX1
Ic6HL/SUT3pMfR+zrXZ2W/jLbvCC7g/ca5T9XZbBhhWARKZAgWvux/9qA5YrN9XT7/Bw1WyeODmK
0vSrhLy5STz/Bn41MhWjxtzf96y4FsPrPp56l6gkbqWepf1wNx+YNVpxM2+DJ6rv1yfqlFYGFUJI
xgSGV3139GXok8Ea+OkPDG3lOagJoSTJY3s2CSbohXTh7H9YZutpu+6KcJYyrOheEVIwnDh4UcxP
cWzDV6AJaeBTJKSbH6zN5y3BesY/j+A/iaiW8ZSWeShPelXF1dpmlIaFeYP6V+G6PTEHTKs0VVVz
uCB4+65gGhpnxyhWXAVSEMwFJ0AG3mih7bYYkWsmpAJoNkZX4w7MmYF47C13sIQQVAveg2QF58bZ
R2fohhGmC4k+l1vYqPs5nHWe0Ap/3385mcAVXm8rv+u5sQIf0hU+qHAdChwG+4E4QpY3VfqYrKPX
YqKH4KTtkl3lsb4OaLWcRheUPDNfn1sS5PoAHKwiPznIrAlflFfbEBjYWRoO1xXRG3Nn9ZPNNbth
XN0NEe2W5T5m7ejCH9QlOdgsgh1dvqBBrt9s5Zdv8IP876DCNC87FeC49dSJPKs3LRWEG1wmEpzJ
ytywjSgMNr+Wd/+rSY6J8nvm3qu71AfSNTArG4+TbG92w3DhA4sKPCd8x0v2SlwAiKPY16WcYXOt
Rja4pMHfqPvp59IpANEhxvkfGed5HtWA1uX9fGnTc0LPKAumPruhb13ATLyP08BbZo6PVS8p21km
wI4aNa/3p7xi0eGJ+EY01QqihNBOkNuos9jkKWLbwOomuRSl9BpeT2SPRNDQ70rivVCXumiw19c9
mn5RwLl3UrZAoeUAGdK3R6hFfPDi1UT7eJ/ngWKVA2vHh2fZ3LSuNJHduh58PrNVutN0V2J7i0NU
tMWYXJW3Mhvm+tpi3Pg78EvCE6O1fgPg/1vo/R1GzXpPh6mfkkXfTNY6oJJkFgUJF+MkDdB4gNOI
TzGLy/jyNdq8zQXHJ7xnyfBUZwCIfvEpZ0wfW47U5cqh5Tb1Bd4DN5uOb/uxEIFA6pugPfqpWKOI
vcKHj0YoR/O4Ffibrc7QOfOw5Kea1oXIajsGKapbS7JOtIcrEsTUpewTv6IqeGu0JLhVbORtg4xL
9hVVkQjjvmGi/4znUcvmvfDcsiZKZbL9ZjVosysRfzQywiJnmll301oVXygtMuRNljC82elASl5h
ddTlVNiTdLekdOc/zQkNLS45daMySzo9Cm2H+jNuyCBmB2+IdFEjAD8/o5FcoyGYJsgITl3fGn0f
R0zJF/Yzr7rrOZvSz7NlZOXR3fxeJOg1nsKbjCGrN6sy9T9tuYGKndipsbd7N4+b3IYYVdNq4Mbi
vXc0iyzul9SdwLpq/2iqN9SqHgTcgD5OyZ46vH3GA0nmWxeTXmzcN5lzut4unwLuaVn7Ve7H9Ojp
vkWfRPUrJneaomM+lwLFNI1zHUZ2l4O0/NCE8Vb9AuRq8mUrSSOJfpVd4XAGt6TPbff7AmMdBQ2R
NKFQfgx4X39Dx8Zt2yI6CorSjrKD5h4eqmDZS4q/yPLdGzv1AxEPoySt87tqUzMGV4QivHTzOp//
hLcnvAqlrGby1cIVATHWr6LpXtLBc/tmPIED+Zl2GmeaYaakjOoWkxsbQHETtk+JNvLTM3nrt2xR
+Mk00VQNhbGtBnfRrzWz/NcTCk4H6VtfEqxh002Jg5MYj/cqywATFGeCLyjL6Ad61/HRTbJCmv7f
JGndhCsK40meWxfLWpzdryes4XT4qGxYv+mRUZYcQxAFGOhg9VkHXcZe8I27d316bjLhhi3s7vqm
jsw2zzjhqoOf7WZHE+nhgGZCaSkd580rpWrANvP1yR2i913Rt5FNmD1BzIhiHFNjvZnHb1wtRXUf
JmFyyel6FL/mSogHXeU43/buGhZ0odCj614BdTpP0yM2iSmKdtK0ROj94VGN4SVYohbctP+TTHvk
MZd39doMDfhTsH9vIMUB7057QRbcJTxA2lw7XefLDbROlEEpjUBPdZb1+Ac36ZRQDIqZiaBWt0DT
KGdl0YNdCriBEcSAcDHbf3xtMiq9g4ojPLhUoOcF+lGfhhH8ZA6aFnZZnExB2Vx7mD8zhocZ30LU
l6J2jMq+i3srV+s/u7W1KGE5JVmNnMm6yQkjbe/vJFZd87NvfiOXiFIL5WkC2bs3nCyRfz4QWiA9
sGAKOGlgIILKeboMi9tmMfsPhSpUAm1RVehxI3aYStygtAWnHDCh4etwHNKabYby1waiPKYW4gw5
3lQdceW8IfzSiRv9Uc4G6ISgji4k8VHfgz9TOjzCP3M4MS2o/GdRKAOI1q+f2TX6HRi2hDCFxyXe
1h/g4NGKB1Hz5mG/pQMUH/EzCil7/X+U8APF3MnW+bbr2/0tDT/jhSt7vFnJ3SrX1jyR0Dcp7Kgk
CV5fgZ7IDXbwOg1WHc7efoVRWIZHaTJWjstOfh/oRbglkfEZFh6sk3Dnr2mQxJ82uEQNNntn64Hh
qvGPHsuPwaaZ+z49Wezjyho7tYETx3MAXHrkKr7CWmQ1GABhxGjSrVZa+W9/5UDgKIT1SqUxZ+ru
BVkiMmwzM7UWRK8Fbr6Ebf4LcPLLvFEqPKhxxLDol0IXNeOOldk2EtgUhfsEZXhO9mbf6XAllqea
vxqHajuCxdmf+Cg2zNQw5yWUaTi25OgcX86vArrCAEeq4VJiIEthb+5sL1LdlP5iNBL+21AWW/o6
cEgCofbksNOouzcT0+77oGtr+45dGLq9WYONKuL0cat6qZOzNqlBnQq4VZ8qcroB6cUuzRnZxQXH
XJIoHMeNihWWbDHt17oRoynj/n8vfdEEXRca+dyXpzIGUGPLdQCkZ+FDu0gS1LvQrGJhaXegJUOF
hGQeki2VOYMa/d8CfSmAi6sXRoKZUxtneOnoT7hOjxDkh3NJO+0l7nnMeBBrMBb+q96+fY15fSbv
GCLcKwLb2Gmh8jWi/GNkbeEx3jAafhfC5gZEx9tstX7NHwrXz5SndULxMiSQA40MMGjUBnLcX+BI
qecCGhpGyUx5s7dgua5suiXRCyzz2ayFYNk8LAWN6kLqtaWk1H0lqgfd4fz2i+2NAlVwoNMTXZYY
uOCGCS2C88eTFYdEM2qHEcRtBN4mGPdHKq0NYD42HPdx+bcf91P1EmgFrwqodHEFWeSnteKnI7Am
xOZet6g3FMuT1jP4eWDyQh0M4DPVy2y9WgFXPULvTrw63Z21zZR4/R+Cw6lIuQAhwZ8L1Suonuv8
/rQqDVSYpaQEhBEU4Hkn5vEZH1QCi4KSQFkH4Wq6NRq0uPDKoHVOUb0tmKQRGYgTN9jPBXcLasnE
xnra/fttvGKB63DabXmcBGOMgRZ1MFiPOFYKzzNeicwL0TQqRhMu5cFibkK4sBeb4nxigqgRYP/J
aViVf+8uIoemjORg5OX94x1myi8zyNQlPd0RoMYtwHOaIAllYH4z1x876l58W1Etxw8jQh5VRbTG
c5LuQxBtBEbxAZBpAGv1ZGfMHVWiMkNlTmJBKEwiaZ/uGpzmZolxLI+GHpz/faK7AvT+L62nJj+1
zHC/oONzDCGzUAjaF884WwEMSbA50HNIwoRXdV8zKDUQ+oI9imK03fhfFvhEPiEKQFndaRjgykdw
aiEw66+0cJ3ps/C046t73krPHxUUGBZoeZPpdMKW8uSd/TcVV9YDi6upTs8qcMKOSl5iZEK3p1N+
4k7CRQAcxPLMHtFsd0yfqhiAPRG2S+57G+X+JeDWhEpWELXYuo5vuRMUb/rpmXIxH0kBfr+ClpQg
q3rnM8jL7ev4YabzSqietRT8/Vu9IALo4J57HlCwFZ0/SkSNcFGWdHsnsPM1Bxy74YWjbBsz0Cyw
rud8GxwPnm0ASwEjHLq/wIaEMyrx4DYrKfAB+Qn/n/cUYqGjEh2n4+UcJQzMewQ6/5FxrC50Q3DY
1isVb2jf8HdxzdITbqC4w5907qpKjQhRL5UdDdc+MJ8B94+7XoC+BW4LBjfiLhfvo0U/SuA/hfOY
MqltIB2NFdESI2yf5cEQGMDSQgR10ipebW5isityiqB5gP7cpfBobt9+OW5qhjdskbhuAAqu4hlu
D+ftv7EFKsT4jPQbArQhjSpQotKAph5QtWT21ly3iUKRxVZT2gXq2HlMKaY9UDXGUEaHBMlaatQZ
F1S+trX2AoxTOAuE+rlbMpH6clZn/Ab75bZYpbHt7qiFlQezRLrZgjhesQtpWsNnUDMkw8VGIPjj
r9TqqI1cnTnBBa3GQszACToMRcUfNcAMnHBHNLa6hIz6qZNwi/2MC/pOftTU8fH1lK6xDAHSf5u7
VIusrIVnh6qRbBcA1cBZWVmkjgtoT7J0azYJs3saGCLhNF6ZvWxGUQUMetNn00WqBxkyUP5V9Zuh
lS1IJDlFyjsDH9x8ZtTIFPBW5B2sZObBq+P39OKTUYzDeemGdSjzpTFAvK2pE7njyl8+9jJiCXFI
7TDt032BY0XO3MJP0FL97ZXqsOoI3FNCBS0oY/6HoX851iqfxKr2cjMca1EBd8FFeYN8ji5wSgDK
KA+c9FkJJyLwOrL0zTnMcOJzcICriS0zfu4qAYbfqluHtNXyIeQYeVolTdW2YFRKFXexcJP9RjZw
QTwKSQehCN2vmeMKwV0y2TJ0t4BX/RUXsEimDNKcu/W5Z2S6qJcwBjeYYZmQdFu38I2xrPlL/G+/
PaN+qQf57pldW7uW7VvT42hbzkkR36OMyUrWPf8WXXivpXLPhxqDXJ2LR7gTMkgy+Y5MiKog3nym
sYHxA0SnPj2SOrKvkjQ7T4Zq6DEEnszNBa4jxX48/AheFmoCnWlLgtdvnVk1nLpG72CDW44xLgu9
kf4coFT9PbFyYGehxDXa0JlWykE11xW2kYQqs+3JB7cFIpVD0tZVniAf2qCSxGwpBoOZ4MZmHKMV
X9azMmcwNyCIQ9+WFr4Q0QCRzYjdgttb5drtz8bxqlsDU9VPHNs9a0lLvD8E7VkoMzJ4VguUleOV
jtsfRLV1Pv01CUsvDg6OqOfkmyNdO56RYyGzLeo8XNqTzCR0IqgYGhWfSE+5UlV5HBfq5Yds7wxr
bBV6jk57MJb2g7OkghkGnhQNKAHmIJOuA4U3jwDy4cx8CZOUTEwnZjQ8frXkHqwiFpuHVz9H1r1q
Jc/twv+SeR+uUCxNQ35aAgct9Oz1tvq5xJPOhmucwrH78uCDUCVuNRX2yTpP87HOTEscQ60N6cTV
lUsqb0D0cZ3NLeBp7mhG5gf9TiCKZz8stO9wGWRd3ZZe67TSGVxkUpniAmoZ/iaT/ffMdPs6fMjQ
x4naOqEdBLj28ekoNZJZ46RzV3gqsWIxn1RK2p3mfWhZFYKamWycG7ZZI5XIdE7s8BoP92NnLNcZ
NgYGSG4kXbmyPxA1zVch5NNqnFx6BeLPP7r4xlxDu1467o+AKBc9wNP86C5wqQjPD4U3FeiXL+Ri
bBvJ/OYnmcq2L6bUbsnihCQn1Ic08e7LixM4GzGjgG7GPWzmy3mhfQ3J4zdqtBnb0AiyXdYwkc04
f5HG5Phny7Sal4novz+0Z4+Pzwzkc4xI8scT3U9K1tFm91JTysc1rel0TORIH8yt/6JAyjGJjvcQ
dC3ct2hbrAZNEBZsKq3cEAvZcT5WY2X83KeX0oQw8THS3MxPfQmIAfLjY/a7f8OpObTd3hb/M7J2
l7Uv0xSmWmNJD2yTs3GznmnbVt7lOlJX4EZv640nuOesYhmO+EW8X2w0kyExTzZTYMrB6VXQtl7V
Z7mc4g4+iwEYtuyJDMXTLtHx6cdLmvoLl33GTx+8pkiIgOa+P3xwwBSFxoRfGV8iVJHcopgghdLY
YwsgStm2thRwN4JZZQ6FSxJiS7cMEg+O+8MhDBy+MR3ORKT9deQWcFLEETBa1n9XZJt/7BS1jCws
g03gkq2C5nP4DVWo+ICaN4tA5HPHcZ/8cGsAdkxys0rHt2v2VxfMWlM2+Qent0GrAg0CZGwztkK5
g/Ive4aiBR/A6X9CX5mHOIIYIEVD6PNKfj5jke3U9FjNVyaRg7gCBwO9cxSj6wSGVVWU5WY3Zcba
W0yuTmtbJ375H/uh7ytHFxJmmpcoaxDFhr42s6/Ya6Tp4cF3rZId1K6J6jar7M05P09TbSMTCcbb
1nWqS4cWaw8YYyzrjJL6uRFzJj3iRd4o28QMD40kZVjtv2To3XDtqsLqq+1zNay0Zveyi8TUljQD
9Jq1cwxeeCkzek5N/IAvNc42KhMqVtjJbn05jQPjYdGDTMoZ3Iy77bbwEr+rd4zHGeG81AHZmrdu
6Kz5B7Mfn9hnHG3VSorH3YQ8QnFCZobIQmCokK89pvuvF9+kwdoqNzbhIcmuEiM5cF3oR+TzdUMj
TlDD4IQoFfdulRbbPwg6UijZcgP/C9Ba7KiNITee9LxqlcTBPO4Ui2Da76w+ULPtFd2D2ivNHMlP
YpuGFYt8wa8BOt3q6kh2AkQqEJIL7DFETPV3LCczXRSIjJlmhMTkyA654woJETgxYfFtWz7UAP/8
7gpwheTO/DygRcTLhNqtMayQHHMYJlLbj4lSSVb4kPN6OPDe3JRxj+lEXa2RUjGNB9Kqoz4l9gLm
QByoGrd2cbJ//skMHzE+RGFlqgIS3vONDHHYwbHzAnDjR3GHtXzYSlrQ5rpNn64LEj0ivs8Uu9e/
rD7uHQR1R3X3ak5vQM9hJhibATJxlsnJDYhqWA41QIKTeGb15QCUHQ04osEETRb6DkEbjdMj/ZcI
ovWvi22tdcGZ2fiZlEBrOWF7ld2NhLoqk5eCH1QiKy3mP4IgBtD4pdp6qOQeupRmvt6CP8XovPbq
klr07zt1RTi0flP8PNmykWO56qRAFBK8tFPogUpMdf5sWi3ZKPEIDZ5244fg71SpiQYbjIMzIsNW
LOWnAPc3FOSeePGY8oitWf4mFVU3AWAr7SiIUqPLt4X63vm6CzKSgh01P7umTFAs8RNWvu/b3YBK
14N8r/K8gV+EYp1yWhf2Frdg7WS8Je4+MWKMVIa936G3waitu0vwSKHvp7+Gnx9LeWaFwuaieDV/
FkjhXtJFnSswveIP7t3zenjJOYHLKv+FCm6m9ghZJlgZ25MRqHritbb1DrOzcXFrQ4LHL5cPRyK8
fqEP5phFuFbijZFsliOaDRrb89WgfD0gEud5QEUohkQVWCsh+zAop+q27wRdxULEZrKSzl+C8Bf2
tjNq6k2zSjMbg2QjxFmt6O6JxoO9fueA+i/myZ6amhRRpk+FlCYAkxHdE+NyQ2zkUjPjyez6xkOh
xoMhve4EwF+QNsWzDN00qGxVu8PQLJZdEUCzlN6v5FCxMBxihezJuLSXFwf8nPGmyPv32wC4VQZ7
2iioqJrEd54T8pUjLr8UHdAoNkNZlhhRb5NaaQGL74d2nCf7RJ1o1jTFddJNgFGIamx/rI8/NBWR
hOGnhVN+0KFpDUbCa16GGdKLwEgrkgkV13qczoMi7taj1FERr6zk0VeiV/Mn/kI+AH8x4f71RCmd
kWYa4HbFy5VVq4of/LkuD0yx3q3UrUuehM+tkGsFhQkrgbGVFASTFp632AyQwjhXau/64s8VHtX1
Oy4MSrFY7RH3DM/jx149zzK2xyzQIRK3dPnv0DftpNfUHkNXz+Clr4ouJ2prR/OKkmA+6ySMQBc5
f6AS/dHuS4wYYmiKD/BFDkKSx6uBQVsD6DuUBDielso7e6BhDx9lEK5pzA67bEzuFKX9zOXDjvQP
11e25h3p1sh81pBqhdm3UkeDq2SY707aFbTSoi2wtoVHCThm3C8lb5EGGj19Jw2FCmVIk+PJJ+RB
MxrmF7MEF3ZQA8+uRo0PfIvqskokPCcPJ7D6z21kmCWA/RvXpHfHxX1qCGDEEXIRzTYyefc9rfQa
d236TGG4Pee1DzMpxMUjLypX9ETrqEPYjvqcAVcPB8FgLBdGFJCAX2r4WwKbI6kjrMFU4NDU4pRy
gbknC5vVkhfuxs44eomRNlJ8wJjvv36XohdUEBjnYL6Z/+Mf1P3fRHDrgDxwpjF9PFD993lfPRaH
0Qkjuv7+QObduNiH/YdEbuy6PljgQeUE01Jrt0+NuCmPQf/qoqH9k/lsB40GHE9veoLlDqYGK6uM
vpJkGy6wTNVPxFZ7fUqahg5o/nDYUdAVz74hTBey3FwbYjpEAAalSqcZ2ey+dYwh67rVX/6aAYR5
ETlzbkwpurd6DqFpA8d3vku7ldgWuKBcCT1niFgy62tw9EomrXcFJrs9zDPFIBIGTIH25AjzzAdi
9Ens0PJKffurQqV0FTMJ7uYFSut5ScVWhpySf9n59a8CN49ua6WDLINqEG8bIcyLTAJyLwtF3d99
jI2ocF3vMeuW/Ed52S+MztcZK7qbYwSTZ2z9THSjjDxnLIkMVFVuxFWpFRrCd3ofHOly7Qr6HP21
zTopLPch7JZ48hOpz0ZbrXzDq9fnHJ2hoOW73Avp0F6+c4PWLsGiLX0eQRH1NESmBnWeXGjvGRJ8
qtnoXdSMel/B5Q3haM0CUkO3XoYR7TyEDMfsOjXqmiSjJe6YcAVA5PRUz7ljYTVzFZcQ1Emyf/WA
7GeMBaKepsW4iHobyCBKQFSy4WIFdF9FanYCMJsupgNpNkk9RJPQaYVkE63LkGfgFFAPkJLdOYI3
Ifi+ufLCWpZpXTBe0SNtGdsfw+6PjlbCtL/wFaXHxxHQu1DkNb4rRq1YHm+/jQvFbo6xXPUe8+gK
D9VFf6N5yWG3uZxAmB9/1TSx0x9ZGtBf6p5M10sHFuTnCUBrNOsHmPoriqi+3zkhXZ23CODXu5+M
/DmgtsdpoVSbp3jgSdsNBrkD2XEoE+vYsg0J/U7w1a9rtg8tw0UWgBRQynOuheHEh8lZKmzXmLOM
hojVcuhvEIBKTus7F/CkBC9nfS7I0QvB0TYG4DQv/gRXaWAHvUC8VFQvP9Bo61XEe193Gg2sFhfY
LNFdfc8U/BBurSgEdOETHU5EUmaR48k6/0TYwInoYrrBDiBprZDjbLo2D+8MiWSD1OBMith9d8qW
1UHTg5lwx+bzZwxJ2AKkgtfjw8jpD5WsRCYsQGqhCklW/wM7kmLBR8WHF5ujWJ01oLXO3WJiaZL9
ke/eca43tPoIgNrh8uQW6b7AgSePUsA8LYte7JT9kzAR6Z5Twr6WSBRzJvFZmmgpwSqTPzYlNSEU
g1wY3bdZc6isa6QVFK9XC0iRXs6oOJl1xqHevHBubT0FAtITYu7A5Z7fuiqYsYkNz5u3gFZyYq3b
rHNNExc8wGw4MWwA0O8oir7AqtmvSmHf/eqUqLS3rZ/G4cpugrBkXT5s0Z9Z0XgQKiDQGEbc62ZB
cjJS2o2qEVwiO+8jl30/Mo2wfXaAbjsr4O6kMqfRht/wouygkjbc87p9vrjuBk4NFQjP7fVVNctf
l/wK+DZsUKjRmvZ+kOdQpTud4poFG+gGvs4lcHe1svCfvePVDTMDeb45pJ+X5z1R9kdV4kjC0OHS
wnUUCsR1d3q7nVR1nO75ErTLDEQBvO4fl3MCaSo5e5u4n/ufiFEG8uCbgOJ33LbuXONteYkweVr8
I3MsxnXWYWHD6igIg6ipTHu2giOardYMxnGXZyH15+yeAqcSTNMQzhkgxFOEUoKUy9A3hUNb6+2d
/4r25Wbi9C7oQOEJCYeXcIcqji1J28EbffAIsMm05ec5x2bkJz1TeEOYIlPTgWQCYLHjWZ9kJd8O
niLZA0p9mK1zpURp+E2jlUWrIRF+DCcvwsl2uKm9jSHxEx9nnigZ8c96Jvb7og0zdtBUTBLScYfD
X0S06vQ+V72xDg9Vuv0EKsBHB/ok/QJuHSKvvQOS7DN5cxLcjd06J/ClVN16tbL94/ZzQnxIKa15
mIuh7WwolnIZy4PehrXRLY7UVYph5K2kYqMhx6q3IPoI5ku0RReMjuyzDZeuqdiKDAbPBIHdCXIH
YfbDz1j5AR/ipnsNrcaaeqBZ/c09NCwZuvR3jHz5g9mwHkQ5ImKfZ/IvKBBiqIVeFFhVKR+v0xaw
phR9ZX60MesertzhXuLalTqrn/stRs3ELN+bYvozAs+ACYqjRRmnOpfLv/1ZyT/ouUi9e67HqkTg
tYkk5K3+gX8o0abw3ozsXEr6CMn4BZ9VIXRgcjp5KuGLZCjF8gGLSU2wnmBECtVuqJI7C88D8jja
yG7boWCpV9FeE8Ep0BHxBUZOdbD4cS0XC8UhdQMfGHNrTJluebir2brU5BxB9gedp/i/qPDt7W9p
EjsRSgVftLrGXWuhTseEhyrS5dPPrbO8NbBlC2c7m53l9IRdrjWoCOE0KfOf4g9di5OkQ4s8hYP3
uvigyr21dlTBwq2d9pDSEjs6QFnRbCfnrCXTDaMT+06OIa7jNkBgrqgVQx+A7sKeyprGAPAG+/r7
uolTIAn31H6gRpvhkQgHeoQB/M6ArEJSZlE2FmiCL6gTprKSumNuxhtWo/pAr/jXTTmAsZFS341m
+IK9X5NkJrVJwCffAjk/6JszaMPXS/L+4EToK7+kFdeDj7qpt8B6zzyXgG6ZBhPNyedgI8lxtXpu
GC3x46C6cZAfhLNEPUKfqoLqlzxKUZDzocGQLhli5uGUA7sA4g2YY8+8Z2OCDeLIAJ6spLlDJe87
RrSzM7Cmj4A3VyYtTrdUpYsXCZRMJdfEH72v5pe95cJbv9kOkCDChBTJswlKFFITXfBnZqy6p13q
UdsWeTnetA1xXEyl9xj3umlRuE39dyc9A5OnDScuHw2bJpnv3ewPhcYO5b+jDOvj6WyAfqbFq3nh
m5cdYotko7VsB6IGDIDB3DL+ZDhNPj2m+A5TS00kZ+C6tY2EODeCIlIerxkS9Ng6TCIfGyqkRQDp
9tr+k0PILUBbMh1wDcIz3l4oEDo0bt8O5YGEdiplQVKZP2q+Gxw/K0TVjPRqOV8isFHtnTgMw3wo
5ItLqnQfdAO7uvQG5IkFwIxyyo2Mbk+ZnjQRYL1i2timtOmfu/CT5vtRtdFogjbXhmyFeEQXu0Bk
lvNn03Em/0G5t/oQ+sVYLfMclcGfA1uBH2YxjLNavhVoUdQCfOdqnZ1g1irsQ6wzY20edPyBFD5o
j7AqUjqHa4LwTKal1d13nzPrecLybVh7hLCMuJ7HJvO8PR6YRMAPbDOMD6Inum3bdMGyyyE8DrQe
wVbTNAL8SOmcOCOQ3A8oEMC6FnrCyPN/ScJC+aP9ByUX0iagQ7VzRWOZwdvOUjDgxwCLe9J6jaoU
OronB6ku2tjDJhMNyTZwwW0160501O2ZdEkf1ydeXuJdpbmgiDuzEpdA3efdIHqelIpihhZa8ceS
Fj72R+VwyPsvAyryWd+H6bF6IjigrFiybq8uI5PN39wr4tW/3CuIbHkeKPNE7jUcP1H0XtgJ4+r4
xEYTITqOs/cJjpw//elTYW46jQbWTfWPBsvhBYyFD8RI0zUMCk73iCsAjhZcHyN4Wi7RlEl+5r9s
czc0NUJL0+brzcVP0tNRe0jp6YaQCFBfBpJrZ5P8QwhLfTx+lVDCqfU7RBzZ+hR5XZ9yAfUFKgyL
pK8bBRMpqUqtKvSvJE7Lg1Vo9QBi3xYfCXKWWiOrxHm8XfDvLtypIGaPBfbWGx51yp3eSoDHLhll
cTRB16gIcKdKjPSUzrFOWFDl2DtIZQdOeg00f9yoUf8mMLIC5Is/IZvwnRt88MNHavdoMsN8OSTM
nCUwe6i14NCoDDZRFOm3U6awk7BjArqTkPsDFBUAxmJ21hL7T9iXa/pdBsp0xl4xL660btF6JYmz
cz8q97nRJy6kwydbD72EL5I3tbr1/uHW183p8sSKhMh2sV9HkGgSfiZDxoYt5fFe4bdDJLHq1B34
dwA7VPnvzyXgZ0TzeYtm71d22gzIfLtZDw3ac8/LGV85k9nVotZ3k+ND+HqyUkW0RIjnb0nEEse+
a/YSNl8HXl0N3qreLPXrfKx89oLtDZDARQ0+W6h9ZD99iTk9uY4+6B0yAeA96nZGANvLUYNeziWP
x9NSDWylPFXgkID+/TEv1daEiR0AxnFaF63sYjvTsE1g/vFhr9f9Rb5Rz30vlr26nE56sXZHRsfm
CKnh8IOfqY3ixQ/+rGEcpHUoWnckIG3/udqXhVCfxYhBLVky0hXHhK2mc/hO2Q4Jgg+zZs31ql0E
hJaH5qbf7S8hdd6LLPHORuaGoGhiRIeKJfFg8qpaKF7sF0B1fBrBa2ufKMaZIVNcqT4QB+OxyWsY
jm8vLlu5uoBDZi7RwSTYmqNKgqq6JACEZ28dB5Q98U98X69ExVf1FpwgGoC/buu5raSbQ5RwOpa4
p0xsGlAc0ZHWDMQmJwpVIdWDPRv5YQ94XxWGSEbm0/rKsC5MEcnIUurPlcD96P4K7cMO+cEq90/8
4hlfA85jlrxvsU09/xyDtJ0K34sDypJzLYiDyCtiSoNNEIywtv6QC8N1Um2F+TrZtb0ma/0d53Ib
5+2EqWGQ+wPPzmPAP07YfqdahFwWk1AqxRZG2AVxTwpkEzKFgmyk9FYWo9ogoAWyNNI1nhhRqjU1
oGCCBev0s2canpIUydtK4aBKZGTDQPjqoM+ym0ZDlRE16k2ycNXTLSppNn/7b2+WrBwy1/QKFBW3
U/xb2NPjYzMFZJHBzHz+Y8N+iiwMoiNTZRkbDxE3NXpWxUBAHy4xis5+Re4idoK8GdQLDe/NqmzR
FlCx7Q4wBw0+0Rn9bzMPmcVtavXhgetVv9T64btXt9sBLTwLRR1HsF4hMspKD3NFrWvhv3oCfmW4
yXQ3sdQuLaSTv9tzJG3/a2/uF4FDNDwZnvoV1U8zyghCy5ht1gyf3HXUykd93TfvCDFiy0LKKhC0
tofdHeylJBZ+7/CrB+Hzf9aoNF1dGqtzlcpaLtVm5xI+qkHtpl4HgueV1elEOaaRyq0JmLEpZJDl
8oMl5lgqjLLtabnWQVl9OJ9PLxHAJqhtEdT6buuwWonth4DTw+Wo3zLC7gcugpNj5H4Gc3dFSoEs
QOUX9iM4V5OcR6vCafKTQytn1bqFy+Ca2iuZCbrSFAynnwmi7sqwRUVOIKyoVOSHj3QiWH3o+2fa
EIWb+GzuW6eE9uPBffwJzJY/FwPdxz6sPMmUuexTt8XiwI2fnThQPGbHI+xFSZybaeJyGmk8q52g
bKxEQnzU/brs9iRLY0MIHRNXwrq1RS6c8vSNMHALR52dmVCV6AKSmzO5ycyERqS/HHi6TPFymTOg
xD8YlK+g8cJwiNIHLirokhFlhOnHHlOmTE5/XgcyUZx/gWKhYidFCKdbhCphRWeBQm0ynyNLtPr/
VuP2IKSWe3gc9mr/mt+HWtZTRtCGnkdnkfiWQ2EXS/YuIhRE1dVkfm5M/QfcWyeUKWN6MrPfws5r
TiCEp2A6D7vZT4VC1yjFfiPkqlGLusRKtgLSTRy9Zn9c8H4mjRIsjto+XWIYasFHwEIUvHGVdLIj
c3wAerfmwjLsj84gsu9qscdpPfMwIqEtyhq8Wq6GyA5TEdggEnMfFX9c621XUZWy5/5Pkw6YkBNi
G0kbemTClLbd/k2jETtXMr/E+yujQpPybEuCkyHqIgdYtcqczViqoBRB+QZnC47n4a4lPTJhtkmL
iMUzFqg/r9NrnwlKCW8DdUfURbL5r/SQuvHikuupont1Ldc3IaO8ltJ0wd0Dqlbasi4FtS/7utpV
xf2vPse6dXu7l9h4Bw7DVFU31EFSnZYGcAV4cOoaiwLOF60EZ6evpkS8mBMKIlCuzWtxrjtjaNai
fVbbgwZycqv3evaLjkIDaMgVDfzn5+kOS2O5o5mpTca2NUjFB5Xfpfa/IOJIBhs92GLuIlbtGv8h
KAuEEj/kbcVna6eH2+lEMQVIQihZyyrnfmJETA4Dq4nGdr8IzA0LqnBdRtUyc2tRtRJkM8ahZM7z
nAsEoCn8j98jRLdPUt18rWU5rh/pJy6VanyDBcyAznVDlN5e8K3w6f4aO7e3BocdpJ2zDpxs41fl
ysEFjKA4Nft5O04pEsGx1eONhO1MJL/Gr5gSWf/IdVijynjWRv4Gr7B1uOrgC/fxWqmJ9fDKOcC7
C7HJXbMEh4dGTvxwPDJ4XocZWg1gL4JVp8GShNuR8C0wddCEJu+/lueGhomRMr/XQwrD1DFvZ9Xk
S9JKs7TcofXyQa3E9i840NjTN9KfT0nGUhuKNXQTTLSevKtv36uQC6GDeCGKPe77etKS6Fd3aaqu
0ww0wtJKBQVfuUzgOMjhnL+pvt/uBWsaAprIsrNjac91OCud9ppBVKHDPDonMsJeCeuBP4iyQ8zm
XYkYMDSu+AtuyYnQUt0U7qOuHfjbCUGWtF8Gy6S8SDm03NP9M98+oLnpxkb3MBN52zM3UWC79/lL
05VLpY9qrBBazcufAbvsM2KaTH2VxAgYJNG9Tc4FRTKOPk8PnmA9QiWbMeG8oSpNChPaTdp+YJHE
15mLOsQCU+8/e7x32agb0kn0llpbKRkV/02uoDlyrSiRMCFhXpjmWzb/L1iE8RfeCAvvJwbuEo5i
mPmJRfTjFS/3xXrQTK+NqB1/pfWKkBurX8pM6o3s2FKqWrslviu/6HMtSpuQ+hXjD3MK+32w+Zr0
mcsSe38dWxMzyCFCX8nWiU7Dkfda3qltnEDT2lwCy38isrv/VLeDDEJU318EfCcoEdfy7J6JtOZo
gW1tbH9EnfG7crHNkottIa9atkrLLNKnNY8j2ha2xjKPNvSqvC0oNPkOevOqiglr33PjdmBnBYZf
nPFc12jjk+RpV6MWbO7Iqv0yF61afnTZudoOoc8tdExNW0Pgo79v53U1Q9qosJyuxkVz/KIgwiT6
bFkMZVpOzvwGZQbTnQzW8XPoWytFmfq50elwJbVF7ZaTfUToPKz3dHpCS9CaNp61NptatVZCMW6D
F7Mh+16OFaVKdauMrDcgRg2YXMC6FIXgtmURXGPOzrHOLsSz29/Seog8CAc27szM+f4aLGAx7JYy
ZT0A3/l5glszoHaFFfZ/HsabQwTWsp1dDKjzZ88QPd/AKCfVKUNqgzGnu6j/RgYWMvEyDyjdZz5Q
U+QawNAn4jZBdPpjsQJiMWZZIm4aWMVFe5Kt+9r1J7TifRVKMiASqFAZez0N7CsBZPP+gEj592j4
NM4yFS1MeLByeJDVFm885OwPjWBeVBfddiJxOuiTZ2uSgB4erI3KBa225kggl8XsDtF4ygGSYKE7
qHnktJY16RSZHUfgbRlvynl70JjTLsoG2Dgtz6Ey/1DhXl8LOurMZNLLQImsscp4OKiC4WG+rmtB
YjCrVvEEYgKLbhXAtvCdX//vlwCyaAafEmHztc/ztUlZ9DylW0BwpbLgJi9q/LWZHLJ26qLlMWos
6dV3Rf2rq2H4pm9MTCmLDXI0w+mLCCG68e3CiOmMH2x07hW/rsriNHEZDRFSq9+x+0Zh7z+9E5O9
GUGVlexlpMyRyZm+/k3i7TLphbvkALIg7PSQvBdIuVIE7ZOdepdPdMV9HrOTDBPNGXsM3H2tWu17
QY+wbYQoFeNwQkvbGGKU9k/BybrZRdrQXms2Pdph0SQWAp4IjC5cLElRlvMzOpmJpMFUJUR56jdJ
7qK+A7vDBSfaMyB4rWb4tr3FLydAfHxqZGNsuSyOdTCyEEtHEVld138pJkguLLj+J3ePwIy3tf58
XdY2F0GjST8JkS7lbfDXx7hac9q6r0YJj31iO/3vAkxi3VnVNIJ9YsqDUd9I9KNGE6sFDS7qa9/C
4NShrz3bSRsQ6kJ3VSYKWcEcCUbOVxDvb9kaQEkPqRBekdhrGcBKZiBUM/iJQ88NlX9kMe/WiWxD
yQfIPkZrgzbp+KVGjh+f2nFr2UtDp/j29qkenjVmd29HxsWiyLc8RyR9A7xyOkA8voMoaZy2wgTE
92jF5oiYe44ngOXYQP2SwV67uttNe+JZH3iHhWYtMq2pb2LZbcrAtutyzvj9gLQppjVQJ1UgrHEe
n7rHJfRBDEthtVF7R0FlknjE4M9DuNfr1r9rJjJAOwD7SNwi7O5AxWWCk/MHmemCJGX74TgMnt/C
6ECkPodIM6DTW0cVra7YKdxzmtouiIImp9Lou9Aaec+lakieYPtr/gVypnGMoQpT1UMz4eBDj69V
cTVfOCr+04F7OyU+bjpEbGtYLDQ/aXzSxOo8jjtC2kSFgJXgFWxhfts1Pz96Ck3rZuKU9bY26wNd
qTfhCXJdt6vxFf97EAZz+9U9/A9t4CuSnJgztHRGWwS+gRDJHnYyv45c+v4Ctq0Oy6CCbFj+VMey
WyxadTIRYJFONTP/NnvIbsO/MFlTn8EIXuXsiSiXVzh63KB72VvYoWsxKrZQTY7dfayObUeYjDXL
tKlyi+w9c80KfbLctwrwy97jKUGqg14/2P7ziMG+ee0SB12qMAH+lwiOL1IQ2rF+EwrtiSFVuZnE
H+LvwwVZS5e95Dh7nbdC2jGbPFoO3EEWwEZSFzABUvbPpZ/dBmhsjU4nMwC3R/rtDSTzro9wvQns
WrRaEsDimfkpq9KgRrBc25Kt3npw25k52HB9WZMy32284bSJx0i5XWW6bfXTuGLjNAA4Uj5llHoH
LJ3Juv/9vlM5tbGzOtbDacwA4qAE7TXRBIco/ikmSHMGTa1GsiArEru2om64dXHCC/JqKmy7kVZz
Obwgj7ccZwxgjfkZwuDAmCcts1FyDgTRYziNaFBaSDehhxnAxybAI4Rxmi/SiUw+yeKASnYSUPzo
j/PkKnpYhEA7x4C+yte+jGb78UsPmYI3JJnCqH2RWoBlhRbGwQHNxh/5jpOjv2WjfL7s81nZejXu
UF1icypKi0R0wOir5jfNAoxQVbZpPuuIgr+xNWU42YEpNX9LysY+5fPXEJsxvWl/a0N2Fcg2WKf+
02jH5O2H5UqiIGUMxv4TbJezwSId8YQ8w/U2FXUkmzucPoCK/NjrrC+zHRKlLeso0PtfxIzF3wMa
fYQKbu3lXFmCdlSj0NRQCLvd4mbipXKVZUAjrJXwlGtx9jE9fx7u1rqnjgw7wwje/mZfCVWuXKn7
vp/TalJNdC+eCt5GBCZsSn/w8L+fFpx6GZvLnbOQxF6m8NN53cHkRhVtMpQA8MZ8XvTJdlmINMc2
DQlYlMF2N3SHRhJVs+NxVu5FmTWG0NI6UKP7Km+v6xfzqIDG/JtXe8qNGCq0u4E6J20cEzNd2RRY
allOjvNuQWRP7hlvit/FKS7zBHX/HC7hJQ0NjDvJAnTUjD9jlPw+8u1wKeckMrXdTMm6YECK8bWa
DS8ofajgkx0ZnVG0FGwLEnhgKAm7bUKS+D3BkdWyScv2ZJkNY2JY/sD5tUVrp9EKSGTFVc1vIK9m
YJxj/ZYeywyGJ3g6jzEc7Wdcu8SY7kplNWj30JAEn3y2hwc6uwW1195Z20KVx63xthP1brlbQdmn
uefrw2V3hS/KjwS8zHWpLiFZx2py9+1JHW+EzEwjceksa6HUIl3C87weQ7MTiWqJUXyAhGEH75jg
BUXRrz/UZOfppXZsZeFdb3jErFwolcXsBskPx3SBbEwdLeA3zBCvKHAm6VnlB/ps8uFbEocOiXdf
xW/BGxSthMUZ8EEjdcdHaYzLn2wWMaBlWb0ON4CTO+CSy6B79rOmWuli9f+fbVnLX6EdwP59XGME
2sPE2Ip8BADp+smq0T50sV1E0Q6BDNIlcjPj7Kp8wUnEKKIS6DoRWaefThd3af2iK58mSIX4Pqxg
jWTeVTxBx9XxMfk9MjZLX8AzVcuglFZC3smQ9KQsEhzeRy87zn9j4PFXKw3uXsyN6XLsq0fo/7dc
EqXpTmOu/9FKT/LJXopKslU5JF/9eoD0V3svgb/TBKQvn7qPckXdI3L7ifAf2ZprN0aplj5IjCw2
/a2+ANUCT0T5Y2dEy4un03wic/eLSqx5auonx7jgA2Ng2z29bb5dgb6dEc5oD1XYY+MGvDXs1gjt
GKbTY96USPFJ5rKmLaCz6F26XP5thv36VD+Jf7h+nsNWIWRvEssBpduuc1SomUvwuxj0J9/d8Glp
52WDB3Exd6mHhKKiKyxYFLhIgm439JXUiwAVD8srlvfV6W3q4cbQ0AYV8k1MEaQPRJR/5PRxfe1V
+lmWv8SSUgMctHosYFk+9vmANtYXEyakbeteLLIPgZGidqhcDuvfDyl/WIwaUAKVG4lISWDgte7M
mVy0sHctPIKOVK1RLxr3q+3VN+IpM82x9d7isK2Wf6toqESwqQzyQXdMjv07i21crEC6JuOK+bI7
b8Gol9ztHclGKo6MCv3oyRSXngNK8AQc2olm9IMEkNAjjS6d3IJn++dXONPobyS/0qYdZ4olWXt5
MC67lxhbrKZPvA4wlvvulRhlJ9GcfS1b2D7zmizsNFASzIL8rVe0xmtTa7k2PQCQ2MkdLXR7IOXg
J3x/j7/wGCt01SanYfzqWgH5v2cE9pFkUw7I6hy3K38B90kk0Rwfiqr9d6mS0YSSEC1xChmajeWE
SQKIkF+vB7QYE2kIaaqAcB2bvgGW8wB6x75ywIn222MlM2cMKMrfZKZjS5zymcnKVlxgQ/U3ROcT
A11fhT807bVbnHinYfliyUEOx0iembyXGd/xSWUGVX9ey1PeD9uMjBTeow9mo+oIa+RReauYeIf8
A4fvoO5J4WscxTSjpuXjVOZNCD9IyMtgKU31u1OS9iPHXySwgkMBg4u3IhCRj/8TGIJjMOZvMLAE
5giBFKcJB32ZnTRFPsfPIzfh+QpT+Ovk2nbwwAnfOrnZZ6jSUbETIdAgXol1H25XZyvv542Une4n
9NAlNQe0mF5rWcqbOnw4yfDHWsHsuuiKccPy0/xrvxASjpFv7O0vdgITGzw7Kf9y3RnDpJw4p2Ld
90XobALEtdH2AmCNYOUg9cn2lZFo9wkqtEiGunvrL1dxCmk+xXNfyZ1tGe1lYRMF+COwD/GUUA+/
nwBNiskDoASvbbrRctlhl2qSpMLIl41aWX+alHv080guS15a0JpSTWDoSzkXF5L4IkX4f4xozPz3
TXZw9XuoO0uqH9k5cin8iUFkfOiNkXk0trhf/87TCuh6KBx6xsOgZXS3SICaowutJy8K8KxvNeBf
WobbthoO4J+pV/HSqmchGsKKphzS343TH043oSQctpydFJ3cVEgIxquCFkJmdYu9OBfd2vQkJ5GG
0guOV5w1+mi/Lu7IuGxelVj5HIM840CRRggPxMgrom+Wq2Pa1jLRcTymgg8lR6iVpwfS/7G1BrRM
z6lL8luqChDepWmIFl/nMmFlig+/luVBILocBXTmDdH3zrVkZCWYA8luJqctNzbkPBNljdxyoPA1
KiRAuSAfP7KGaslku4IJsLmfLYYedSvzk35FFLt+2pKc06/4rzoQAWXC9ke0XSbyOgZINwJN7ukN
2iq9EALTnoxWUULOlgTWuKVy7zgSDJ24Ga9XHSV100c4A4suDI7K6tcVQRmKHdQOHnrdIApuYcXZ
9EdY1xxrgiw+HnEnfpU3BPa1Lh8LGWR/AKzSkFuEQgpFHKCc2tp8Ibi6K4WAqUyegQMOTzL/NbTN
YbvkijaE93vnt0GBLKS8+hPbCS6AVBBwAigG1pbQHP4oLOU6dYNXpy4eyrksBIT7FvUuHMMEGPCq
2EalfooIb/DTFPWRneEAtqKFJpOwyZ49sq/xihCx9MHXVOqK4c/reK2ep6iZIAn/aJ7wRNb63U95
cdjybBviH3kOmPUJEdTN7qbPqh18RBFp7cZTvMx23E5kJw0zuVbHef+IR1WjP+G6KP8gac2Nj5Bm
qNx6sc5/itje+XInGGHd1Zxd0e96c6+s82hiYfHW71SjeE3HHblasamWbybnIkgvWc/lRRbvPziG
9V+UhslbwHBEEZDkfERhwe23r7cemCWe13rflhWtpi3uoNnjyycu5XhhOJ3oA7CqU9H2SBCGu33B
F0UFWUFr9uCFUNo6Nr2opqPKCotc7PpSX2DkN9r7fIZwRdooiKqKZQ83LkxgmIErN8dy+E0XGbPn
19F68abcHrcBS5Grgo+3vkMH2g0TQdV3xVSKbKKwLI5vvJsx9An2e1GkZjGOGKfcf4aCZt2efV4T
ls/qk91oielOoZDs35BhB7jXy9vL68wr2tLxueglIDok0p6u86xHbVZPm7PLHyvY1BtvUg5OEvb+
woioa8kUBbYG/uNuw6eCrmehKAikdqzCGgGM+hlUSw0Q4pBmBHaDDO6rVJFMtHCWD2pAPahpFPUs
/1bsmZsQ0SAaSBxR+AnHnj0qtw94e1PNXVaDqVo+nUDt6xT285Oe2qV3mdTBvLLaVXtnrvEbMDup
4DtkSB4uNFYmRaQv1mag/P5A9+oEKb3/818xDw7MFJgVSXR3DtUBPKNaqTBQke042m2sZlfiAwr8
JkMBl/hOnby0Zf0GepiV8l0cRL6vNsd4vz+4C1Qk6fgqUdqspy/01KXv0bZHYPCa2bi+fAJEwDoC
akuGyCiB+/iQPFR5HR/HmRBAWb9Id5yqrmTyyKEDg9AAivBfc4CFpFx8xN+XRdyPQWhUJWeOEXjP
BjdJ/QJtJLHOdbhz5FMDtygUUYniRZs84lEM2FX3tcTRIDUCAwGMKgej359vca01Ekde6rzPBYFw
lQcAEtiht/G+0S+K7UDUf/7ss/Czgd8c7oZtcwKQ6SIrogIrKf/gqhjt/ou3k5tYNXE0QhAw+Bxs
2LMxvog5i2iEZSR+sDqxhpORdpHdPTNmQIthOSI7jUYUiRWZ2Nrmf7HExpg/1nBYEn7dehAqmqGd
T8WBWiDxuJkbuEFryRMtRmpBdeEmydwmugSGYgJ0oIJvcdhpd8ikQS1HmaihsN6fATvX6yNVVo1o
2AOKW10HB+gSet3Msc/L6PTPoNcYbUQ2n5FMXuP2bvyuIezoMiqDNoNc3mZNbAn3LbQs/2q9uYX/
H6soK8AYxR70VR4Chkp2DdkScpKfzG/nlTvLdz2AIM+y9XjcJfv+y9iNk8IX9Do7hOt3wPiQ6AD2
Ihy7HHhn69cMh346Exd4tN0ZbgvYUDkyWjHSUc/rOt7shldwl3vl1YN9Tg5+b7jG8YGzREmHOaU7
CBU+S7LZjp20mLkFPXOL2g10+tE19kqMKbLPT4X8BgJNX6MZ2oT1wFHH7Y1r+8LmsTQgtBdCbm2p
G2rH+K2rLgn9fJ4u8XWFD0kI1WQ+0b463TwCEiZFRRVkqVeBnUh131TCMRAmVKoTiP9Dfo9HEtBC
pGdmNdF0NZd1e9bcMo5/eajoHzbJtXa62jMd7T/dunzYx+3qtvQeE2Bk0Xt3PBj1Hm5r2+oUyyPW
Bj1ZBQb3Qubl0Dmqq3iWcKipxanonvFwZKVjsfFiI2iaWmc1peVrVY2YyXse9gB1/bgMKW/jju27
JDeHdFU1DMxJCmc2d/t4EurP8JbASaMJzqnXQpUs1fZctJGS9kXxBJ3R3ULbbdt8poNtlBSKJuLW
Lsi+1McyEF7thIT/hDFHRcpvA0iiyurerE54+OeOSRxMFGDPNnPZhO0tftMaGC2OoW9d18K+u2UP
fVI6UDMy+g2U5zCCdhcAXf9XT9Zuq7niIv4rYN/Y/XyF8W/hgmNvgcX8HlhPOu2M5uB8xhIwn5pZ
/F8Jwzck5fbLYYC5Dqlp1FPpwnmWrLki+zMk6JoWby+2cGiZFxv0SLAST7SzouaEZ+mdXaMau/0F
EOTbvdfG3AV5DhLbRKPOTouR3jFPlkkxTEwNQ539hp5my/WSKhuo+82UbApgVTOX+INlk7MqqTyI
5+Bfg/TyNEIbHxHq/sfgtgI+vR5OgkDpyoFb5zkb8p7FizaYLZ0uSWgEYRTUmfZ4GVn7bd3lC1dW
zPSrK6fC1PRfKJ2YTa2IkjN+UU//C1SxovI/odBUVF5oTiQfXMf558PRqvumqJ7QT9gtV4RWc69I
GtIxJy8R+HW5Yq90fcwGZY2aOK+Ug0mWiZCQ4TxnB/i7G9LiqOEQZ7iCIyxm8Ar0n5lZu+dknohj
l4HKr7AmyAh2hIX2xtyEtG1bo9HTQMKB5OjMGshCYXAx1rl7+xvTP9B4w3B8WpBWBkY70NYmJVMO
kPWvwXGNfr2dV+LFXT5lnn13XaA7FEDxPhaDDEpIwV/gQ0N0KdW5ODRYUKIcZjzJnYkmVs/uDaad
2wEqfwPYLQJuzjn2NNZ4K8N7f86V0nVz6i11RHvWQyH5y9m5HJ0lO0K/Rl/MQLJmmfLnQV6GudPf
adlflbwl0nmB64mxP4VnotVYhTYBNht2/5L1RlTMiwBCCpia/+ij7Tz6WOI9Ad8CcUjtZPDYpT91
SrmH9Z7EtcHnkjwsowaUMWYrfI0Kd9c7KsBPrw0mc4+xOesffobLrQitHeq53mhVss8PmVuBPpk0
rrPj0KlO6GpJg+KozOvMnXzsuXP/y1/e1TIrWsqQLXGutT+JAZPkCbOI6U+tWFoSf1Pe0tfasoEb
+WggsnMhullElRXtbOUs8+rAN90qdSLVrW7DnPn9winAS4qHe0I19Bi2I4/gQYS9+2YzLgkasgRE
dTeJibSjfIUQZVkKKUdBwt/hYxRz4xDn1MXtxOrLtcmnBOOiKARmLEwgo7HhX/kJWd/h0g5rZWcp
EneUwRdcRhmfEogqrpI62EOd+akYsnmFAhdUsMCTft1VK1FTs1kvB9e+CXe5KjA7ix2i0gkzL01V
0rE1jcN6IQVkeHsBmty4iagIA/opF1miwKPL9xWY5xvNQfL5AYzfLszDW3OX1Cp8gFgh2Kkm1GLL
6m5xD4GMn02mjQcLP/rxNCtNoTClWLWj+HsUoDkKrf5BD3yVX0lXaRqsRpqcHCHdHUrp6gDZorzI
YDHO8pSeLdmVaKHaJF8fnVZg2usFeW06FkWF6lZdqH/q003d0l+K7BU4bIBb8cWRszKOlkzE8TFT
xbTlNJTI0Px1XgFIfijqDb57WuCuJyb4ap37GsXPzi50qto/eklMgp38gB33aJIOsDYKwi3g/YJT
IjjLtcA5A5otC+In5MULGdsOcXmE5UKpbCYZBxHFqizIcQRYyxjMus9Vo7r6y+smHtY5ilMTUOuZ
zkZiKBgy8wZJvrnzRpNqOl1AvXJJgKqOoDPGDq/wsWULDn7qW+pX9sFkSm7STxRa4TzPTqTCahmg
3jbLJcEzeblm6+6fl4l5gS4Uy1yyiT+bdHzegjfStd7qFj8KqvXNJHS1tz3fVToK+Rlaw0V8zg5g
026m4jkTgXxtGRjkUnacjPC2YadcvQNPN7n2yP+v765vB8G9M0rRwuEAWE/iJkWd6BWhacH7NvHi
RTu/6697kL4p6STpJnNggLHYpgpvgAEU3jIveCo6Cp2lOgAHBLMgpdMtgMWkcDWNw/0hmYxuHs+d
wsirZE5qkmZTrwsq6xfnHbjuqX34KsFZq4mJ7EkFC8k+Ev1mSy4TOq4/+WBC/yq29E/DNZJHCDfK
xva/VRPNRvN67iX1MhoOntrWMFbLI9bFhAVpxRUFYaPKrSZUrQUKrPQ70XMkor6j/xEsjAvXLoHn
NdDUoewRmkO7SGr2uKQlGNcWsbLgkqKJsckQ4jmqmyO41wAU6qLJkRpU2f+XJfakcWg56geOX5nb
xpxhZr1zTgH7I7wSGB4kJQFzVsXlpaXLogo3Sz/1Zhof+a4RSbsE5+wZY/32HGKgSsAFNfEIsTkU
R6mZHAa0mn1bE104tH/5sevr05jqYEswwL7xvXXV82Tf3Q1lkb/dVfnc8L8k4BO/ddyjpKQ9luDI
/9RwGeyeokPBcgsfhdTpBmNtFaLwM3Vb7dHgRXWEQoQpp5boh9l0auu9Tb8eohLE4tv7+Q6qtbl6
AOo9HBTie3RpfzJdKe6VwNFnX3UXhZYNpFeQWhoNpPo4101nY1ZKniTkalErmgWeKOaHDtXt0ewP
20BGYAxev66U/f5kNOFnK7ao6sCRc7TwUgRaH7uAJhTp0VSfaeKanbOMBrTnjcljgJHxcDOLzSSG
ifRFXSmhlIHbVSBjDR4TMx7QxWQc+DG1a9//D26i9QdgEZLV1XPDjCapIjI51yFqT64bdF1juwr6
Krw8ltXh4/cWbIlhUXPQKREdIqohGCS45vpS00p5YpGbBDm5Q+3pMuaAxWRrJhM200AykpC0fMwy
gF94qquZ5NCZJp1iS1JNFENGSHBYliMNdj86uoFTRpr+/qAZr6j3sci7xBf1zpCHWqPO0gC7rflM
ROeUevsL5Uvq9w8j5KT8kObUa5rK+SOFvkrQRGpVM7NC5cYfG2snLXJNNWP6csT+3xXBiIde+JJC
8aFZkgjAan3vg6QW6wTl2Ixtay+TYJJ6e//VmOGbmoF5IKW/D0knm/mpHPZOoA3LPqBc3PXrkJ25
ZyU0lbAUA1/MYg1QbY+9+8zNtFduWQmPgxyqjlJmV/UCKDFmzv4NlFtouktqLPOfgzyFnInSIosD
lWJ8POcazEG8wAyCbYsTGGKJB944AOwIr+MWBYOkOjQNU2ELqh+YjIILvfnINi+YoWZqMY63/BQO
ER7Gtazxj1XPISzTi9iJUuChsTsrhzPjfNNlOzDu8MEWAMNkBLv419XTAuLGFwbvIi7ja81BqhYB
Uz8+QUfqqkqQdphTiK9Q16gtoHeQyyeFSjX+2cuYVhS2yfnPfomQZJcG6Db+I1FT0IlYlEjBkudx
2MNK969bbqcv6anKP5XBmCK6hHwowpYt/98XZZWl7517rwM0p3ZEXDMgul/0mTcAPZT/dIT+AKul
8dzaw19FgnWPkV2rHtddQ6J4vh1pPIuI9u5vb5c0d3IGEMMNKBju8FJ78L1502cJWM++Rr1NFjvh
IzesM0IHgxZTLKYurFMkCWxAQmYRNZ3eM2cQai7dtxOeH6Eq/qwiY4ymX0TcwY5m9Iz7otgLw68b
W+p2+wU6Eg18mVMnw4cr9+guxtU0frBAsfVLNvYLFp3Yf3kYBdOCVC2ZNFmuOTYGZiBryrUS3Jab
STfQ2v+NV1blpIvZPdAPCwBK3nZTfjnbTpdtPtXaA9EqIItiidmCFxEc4yzMsHrSEvDUEse61iZ5
aUhqpP9bMhkWnX3sPGBvvCZ5I1S01xtpCuPEz/EQ59c7cTmtgRNDT7tzc3QR+IRFmd7YX+4gDfze
8PF4HVjzn1QxmFDgucVMaWO0j1lPXOIi0fTAdcdPZJpx0LwkSovrhXzLQ8+M+M63ycY0daLNSzhj
cVazgnFaKBALivRzAaui/9q97azDPS82rmLWN11XpoDdT2Zbbskj1XZxHvkGp0izFlnmjvqGwnsy
k1zQiLhxmKqBi7/m2F8n/n5ajLQIOnvVmw9Ez4k5ZmQ0HEqQodl0ZwsciElq0xmWuqzUzK53vi4C
Hydpk2SpcgzIEDM1UM39Yc76jXe8fSlxpXtGYOp/7FQnKg/tMGMYPsI1t4K5Ze5QVHHfyseesygu
r5Fm29LMcmHUQ2XGkU1PWvKJCx/PtnJoCmnyT0cv/4Feaw4TD/NDU9ck2rFN9TToLDxF7uoFeXUm
rAOU5qWgH8vqQMt6+wOpGV8nyhU2QbXJnemGH6LhIdWCX9xHxpNdNbvcqg3LCzWy94AgoVe2Ggsl
0SdhMVPOKAitnAnVA+OeMhFmayOROs1ps0mMbzuO3Nt65UN/bTPYKYrQJj3tNx8dsejkP3bgs1Dk
3MMJygifIL8K7GBX1wAVGf51XZYkVcUua4of+b2TmgaMYX9I6fNRzDH4FV4EBNxUkeT8Qreb8H9l
UUwlTkgM9GxXvCucIvlUvKuycP5tCaKRU7QdjziT2bMlaq8gSIsJYMxO823W62BPCr7XRF+qVLV8
o7axD7uZF3WcH5AP2IfSMr3nPEiN6s/21LibJcpkXZBSd3Y8DEUdVOI4XFQBt92wG7i7tNJHLAxK
dkzxoaOal7F4N03O4PV0A/6AQUU0ZwxvEPp/7psxLGDCbVvrd1LyBYdSGdmfteM7Xrzn5lqUPfl9
SfUbPhbGeUU8NOxXHB9Oto1w9IkBRCzIkBBnD06HYgaVr/8d+cODsVXwZf+BbsrqrpzaSjC8Npeh
ECGQo/4sitDjosDpQcOKMPz8jW2jdXGO2s28oqSWkweRz6n6HDIyXWYp28zwuFzz3nGiuzeK+I3z
hjfQ+EmT8+CuzxP7+8/MtLlV4ejjcPCFsFoBQPbQFMsy6O6Lp4QxPRn1OhLn2qQhVX3V9Lns53cy
JmHmXz7kPdjZaAzMX/o7KZN+4GLgq1MYpajZ9Cw96tWVzoJC5YpvuhOSga2UC+X/Ic+Dt9Ogx2Tz
Z6JHVRQ235yUSrwkiamJRW1fxrXr85tfuwU5rGIJ/AUY/dI8Wm6TSrH8FJTmOG2yaUflrRmRcRKh
AON68y6gNjA+kmUx2OVC8OC11kG1RYfZPvD297v2LAr1Y3lVqC2AqJUY6IShhxOipv8+bjpZoVcq
aQDjuvk1H+erebj1MlS2g9gY8KsjiJUDbg/fUnKM7RbZwOO8RplVdW6KiZzRBSJZXDT25Tn6hW0C
fS6GA//UiTQ6Cm8M/WzD+/IEeuhZmzgYJ38hF0ekXCERtqW2P7UlQPnQ31cETe7FlIw//F3NRq/x
s1eiQQoNeFh52MdGKdVrAqgkraTIjlZLWdVmUMBsGEqRZXFXkfOViH01P+Y1mcx8/DKPukNVhJ6g
MY6qCWMwVlnCAWrz8naPNk7Jn9zkqj8GYlSbQjwuitdqe3u5YNqZuVkviB1hr2Em4IzOYSPAbCoF
B6VEMt85bOHOh/gFztm8et9JFOz7lvR9LL7MNGsZVGtUdpHol4bKTDPXRn0j95oSMURL1jSqYIac
LAF8/3czFzz0gsoIV96bjNXETPXI0kd2cBSdJfyPY9a8EBzuuvNSlBKKEIA0buUHx6UO96mNajJt
ER4hAezNE5f+caPsCvvxbT9tMhkfFKtLCLM4NNVJU941bsTjL5i5SZb3tvxv1TGIHBdPrtmdtIe6
rHDCURgdq9T+pcfpHP6ZQ19EMGhun2H3S3w7gPQ7zfIYl8+ewBGsMX7TjguFIRpA5Et519z5c1OH
d9ifN0a9fLntcco6nZu8QC5oHrnKnO0/UyBn/W+BbZBPSFAt0wugopP381f1lN1BiYEwZd+9ZzCP
yO782cR+R8rOxVPaQ9HsRRRh7VZ3MTF0UcMMYfiQJ6FYdWy4J3MBT0+fu1RF4fnzp2IdvQun8QC+
cllaoGFBvC119QQTbMClJt/6hpQjw1p/6lBpFbCKRwUeklcFsAafenlsb4m1W6lW1AzDu89G8ir0
sgK/N+ifHgHm1wSY62Op6dJL+agBrnVeMdzPZhoYtLZQ9NvW31VZw6g3NDltKb7mX5Hr6JzspRSA
2r6YMIFpTtJMb2agFjJdz/Ei+WirKvvasuCnS0tgRoNVfnm3V1PzIdYIuYa/QKvvn+tzVEfoe2Hh
a7AjNjzMCNI7mH9La4JsdponDKfc1F+rtVDo/pPrDOZWUBA5bhw7t6FJrtQryD7MyJmSu+2kgqtb
g7L8BcH6CEQToN54O/HnSmSGFTKokpXCyo0BFGCoB+66JutOL6pAhL89C+vKN2L7gw37OW/5Q0F6
UVURWryzmerZHKUDEWv869zK2YY7Ptt15+igkuN60hHs8bl+AZEygoDMr/r7vr3J+xWtNorus8Lp
iOJSCDf3fzlNTdHL6ayesVPLofNz0RATijyR3GmmzykEkztD2p/mqxnSqMgoBwQm1zNp9kolVd+q
AefAF/5Y2x4Ou96zKGwOD+RskX1r8sMBNaPx1/Dp5+KERBZNqibvkXxdM3yj4fiSpDCzeSBQdbqj
H79LJXcQ5dOn4hvg3wPI2A0LKd3T8yEM52JQ2XgSpC6YT0nIBishBSAP3AVaFf12d7pPh59qEynt
OTCDiqQrlkAOBz6Bsq7vBJCACdPKBzasvIV2BpsxZs/Q1ExbKYYqW9bZyP4Tmv8/AYEVzpPpFF8r
Ai4y3nehkeKJvrR8MTTGrxxfM29Pvyg3qYPn2HZg5xHulV5uUYqhhi91B/MiA1Np4Sz5xyjQO79L
IJXWlfvuRv7PkH0WbmuqOLtLyfDCwGchfozyUwS869NL6BpwGUCsgmRS7qJrS1Ozp6kQClnvUkhf
danu+mWi4S9KhOBnIhVZZ0X8HunFhW/X5BnW1jPAT9Ou+0LcF3pXDaMkTv3QN8DpoGObesMzUkpr
ilvEOY2KK1R3JvuMULHksg+TKxGTQMSOtVCro1+UGSdU5JT3rVevoI1nRmNjQKH5JYFe0GngDQo5
BUYCOADkuah5SSMLoZzNpaxnUygadf6ViQpMt/soAap/2QH7978o52HDU8js8EW3QTO9n7tkOEaY
It/VAhH8XeFG/aThgYEhjOz2DL5C82EQUArXKaBNQCmmVzHv1xgI1Ck7Xl52sDP0GMcIAsQ6Ga3v
3gqsJP+brT6zUQZsEGrdhwKcfjsgd384Rbcgsyj5rNKV1zL7aGT96O4/NQybgbvT4wc+py42Y1g6
s3ueGW35KiR5ta04K9zh/4BDyULcR4JbzfBsg/N7OsNJqUFa+vFYkJypyVcDZxm/ZFXtfTeTRHf4
5a9VQJOQXP4feaY8FDlaYx8HG5LiLAnZ6cBUfefkP0i8EkMyJx11pDw4fpNrQbD/exrjMiX8V2Ky
D+4odQ/RU4E6LJK/GgJtkeUmGVgpY8xBskTnXGdaalBJOad+4M1M0jettipya7bJpvBPk40GG34s
Eptus7K9gu8CF+31yYji1zBereXDeGhqQ3reNL5o+wOTbVwmWBWp7XtVDt530O+caQtz6brNFp0A
b9dJTkUv8bnh18Z0Vkr1WglpTueAiyS6RKdN7DLPkn2hAKEXsWqhj3aVxtWVPkWZgQUVYI3eeyeM
5UXSnmTF5i9wk17QlUr1jtiLOx0lcnQbva5GcKKsL3KcrZu8T4MG3GyyP5Lj/TV8gvwUM9LGCnUK
CL0UTbUDxEZKSNkQM5+yYMEswFhSE/Uo2CJ/ejQ1PZlai7RGxxbLfIoRn7wji9Lnd9mpGqeAaBI1
Yab4KSq2dXIuELsWJLzBZA7Uv7ZSNg7rmZMujZgtSOLIADjVMIXFEO/S3Ny6PcX8+F7Qnm9M9mSW
Y3Pq4iRdYOcZ/Z5ykvozMW0c4emPVyMBoRmC1ptaOa96xVMLFqUJQ2FpJxAovi1JJJifP6Jmc2UQ
oIUXakEbn6BmGNxFL1Hc/Oav6vOjyVapcQd2iZ5o3OEgTiUlA4k+bPY4+LTDXdTpATabWK1+E1qs
sGIUed4XzypmksCjaud5bfIEJSTEcOrvRz2PoxCkD7X8Wmic05sVPQXiDsTctmLtwILGSv5E8psd
uYHwww0Qek6IEauLNq7/zn0kg1fzAsx/6NWoDQ/FTgSARlP97KziB9i40Tg+bEehcvQ0J+X6BZoD
Fhp5/ipUOMIOEA85SwjWksS5dxVah8vXRrP8ikje4RuqjCb1T+GdBM9cAyWQibnBTRuJrts7pP2s
lPNG34Xe973cJqEiR0DjUEK0AFmhEOr5m0OxscOiFllDxoAc4mUm0N+n7s/aGFIjGkMIKlIg2bPz
J3Qcy9+6yqHF0FBWOqUglCetarLtCWNvL8dnyKdkxgO1sPNVHB9Ga/LzBAK48kGfD+ecxjbvkmcE
14A/hFO+piPdB2GlyalCZn5gIdqdxO7z7neEW4vuNKc62N8+6jsRxq7QbGLLaTNSIz0ngIP3yifC
5j2K5y7eH04d5E+k+XmmC3AtNaE0+9otkEUR0oY1MaM36ZosSl94p8cyy/JAo6hrCBeoa+5yYm1V
oS9rYJ/Xy7jc1P8G/jR5bQYPWen0ANUpYe9EOseEsV37Ta0cV5KIqvQyX6dmeIArA0+qKI/ccg/j
j2UOuHGKeWsv4i6wlOYs/0BbhOkbPYAGnHCqB1viq2LYOWDjHFp4y7CqK6/e8oKVCNzBo/5omHDY
Q00TdnPe01PUBpKGGaLA3gY8nuO+r0oB51OnU9JgZgteAaJlC5D/wqhbLUqgX+vG6pYEIliAkFXT
bcG/I236SBQ9csDt9ltZBbVan8u/fDXP3V6MHtookWFmIiLoCXPKQ0qZGOAn1RQ4wUghTNwTMCmH
pPXBdYhLeujJeyUVY/di+1vwFonZIps5ptEtrCLYUVFB0AyG6gc4GPd4upiMMjjBe9aT4LcTMB7y
sW9H52eUu2Txm5KFYW8Jh2Lj7bArD1LFRgM+hTPA512/ThawNsGGU7hQibY8U5++izkr+WLHf7km
AQBvIdtJfiglBDTs//sAsQv9Q4JbCpPjmr4E3AgKMFUApzvjZ9yAdmTbJIygWQQjdC8Yh9UIdto0
AeqBzpTmsFTsQn0HvrcqO/K3e6UtUbhb29X0HG7XIk0qZepCIkIbgDmtbErH39ZvHwiBFd7XMAgW
rfs3f1b4plpD+LN8DZPALN+KhFjGmHPFbfTWhBb4sYfDVquHvdeJbZDe2JHXdb1oJf8y1lVeavcw
vJOokfjwyvfQxRlVe6R331Du6gaGCr3egDw5cNEzolJEL6Xm9nUNj6ob5cWk8dYx4c/uTkeynBe5
Zf4NIDJw85wzmRPoOSH5qlAvkzP2lcMNC0ObnHE+N3I3apKY/WT28rw21ZpwN2nbhS4dtG9c0zJj
N5QD/3rgIMBaVO/VYFlps8VVbBigGKGmnowBaoKpjF/pkf5rAaT986yROtL6IXfN+vK99XhY8E8z
o2K9WNcGEp5FIhsJFSekcy3m6QblVxzJd5MLHbcD2tiWaPN/5fvJeorvXxAPi+tz2/kSgo0C16/N
UCIJHza2OlSSHhiKK1HmY2LvZX/NfKTw2vUPKC/l5Cykh2D+LJnrjPJebxON9v64jPaC6BK+TqLo
/jp3QNpBwo6iW/QO0eLos8QuYJNhhd8AveteB/qPBT7Ht9QSgRCJAU87RVFVuhY+z28qlh8RKDqz
eMdH3gWf5f5BcEaBvFhvQP2T6On+N8K07B6NeIeVCKf895pZPBL1rVAPzKnhj9fvi4xQuTFRutU4
GY6jZeyBdzqNizdeUQIH9VagSxbFL8YSIry6F6xCIkHDYFibDdQm2SBHfP37YPRdJGnlWMWDqhWm
IEBe2bP8hhdKTs2LMaWm5jvFYoJzL2J4hCd233Ml3wO7TDcF8S/RniKpL8fPWenIdQjwBrd4MWSc
jr+9sjuCVnNKZPN9Azr4+zi4Nzwmb/rLtlWA9IZSiYsNGdPAnbfJXlAAhM1HUPIS4z6BjbqL5/RC
V5VQcXnp6tyccK+zpz+DJsxllyR+cqpDbgDOpGjAnELWPvk5igW4yHYM6Fb8/d7QAC4ZgyYQaxqX
bR8rbZdttfFllWLPfMWSe0YP/h82hWsXLJCIS142Kzlj9sjzoqmSyEgee4PVigtBuuV/sWBfCT0R
S5s4S3uprPd+NAiHcNyy+7DDGsM7m0768GUr7fnSrsQBq5sALNqijRptj2EFNxEz0wInKB21ebuy
n1Ub9XP/VAUSF2uOfHRuie9/rUT+nUQ0ZguaB4dNxT3osIJfcYgvoLpRBWibcmIIl1l9f9IvJf3b
h9qJ3TAUN3LaeiZVPArkR9zmPjhPpw0fjXo0X47SSKvPqrzCyEk/Dn1Z0B0l1qilvuDAVqlapFuj
Zy7rG8kxJ+bcBvNcmYklQfegcDmZhQQAxGonG3f4zSVNhFNJu9ZDqYYyuB6YBfKxptq8et3i8+4n
NAilaZtPABAtMlEDHsbjWnqBRXYtAni7O+hIGwPGK814sA8xcBBViSl4B7mPWyz7LHEmAVUSlDeM
ezXNhM0wFMQv0CWAjVCkqjoqJ8wQhD1sq4wcbDS6AterfRqPdTeu5upF+8VIiJHB+ijHSY6q4R47
rCj60vNDaTWcniNGjRBOGQqftFYmieJzHv0wcXW8RiVcM2zonQ93akhQBck6H1JXDZo1NvcXzQ41
zvScdD6WP2Qr8FWHlgD/YfH9iRQ9wzpU3DLGTUn3RKcUvhfyVJS1nlfq9HAXVYSS5B4iVV/ZnM5k
zXxEgX/LGXD6z0oXyiFeGGwBWq+oTzDNYle9K78YdCVGy7+abdcCgRJe48nFjyZw+UczO46TELxo
GOvqO9yVvJG8pSBQDfAF1dJjFLZl7d3TdgxeG7YQ2O+auGuPpit40UsFdv8JjNXhXdjZXMczj/AN
25UbVsnUy1/Cnsog/bO5hs9VRWPBnEeHiurUsfE3TyWncqO/f2EuHzB/Yt0LSFVBwQ3BdGGx41E7
QSGiBqViYRwq1vFHnb5ROkETvc3K0nyDsbQ/OeWcrSU0amzxrc5Zv1xFM47DdkTGKN3Tbzx4Oipw
vtJZt7pRed9r2vMBy5OF9vVsmUa7ZLVFg13c5sEa7pf1EYM6iXOS2Si7VCV/fXxYQ7Cvl0r3tzaw
E5S0FFwA4JP5TfJP5rKlAOe1I8oIAORfdj7Nx5U8QyRLzIzRu8xU0poLOqUAiERf0ewM3Nn4KDZi
fRfhMYyGtdy1yZYwX9g28CHjbxnBsusS73olJGzm9DMhhGRt+IrW6ZPtR/++T3+VFiDVk1/HH1oT
4S0thVHqTwwIzjTuF54dIuSegn8gvrIhIHkXT1HaUPlHHk/xkvyRH+GXB3Dd8bAnnKnLO98a8Z5W
4vgOJLn7B4Yn3LBAvnAoAQI0D15NwxhZzqHeS6Ud4EsccB3zqYd90Jhk1lm+/rKvQUhl9mm7g6B2
jxxp3Dgou0lRdeb9iID5OB5eRvLfruvpTeJ3HjcXCKkn0PYEXCskon/kwZHUehomMpuAzYPf2Igs
RZ0Zsn0CRC+YYNNfZnc0p9zzHNrVWbcxOqjDYIhIIosSof8eZ29xf8x3LLcdZHnQteZ3ECcsDRTt
dlIkQlaedEIZRYreTleu3sWVIabGLQcmLHsaDctyNwUuMZaNcZcQxVRNVd56Oct14t5xECQ2hn0T
nh4ifw7djcvrp1fO2PxEcGcPtJEbtuA8wrjJYOomtAVRVNp5KRBUadIgbwhJuqD/FXZCpgIqhU1I
EAn6Gn6zIAc1kYl/jNn86MJQ+Mg8Zv95EaI8jMXc1+M3LNEw+RNUEeW8EQygRSjc7bAKj9w2KpKP
PdoeC1ZwhEbiUw1OQAFG3nat2dDNKQhSGRa2e+9isr2CmuzW86rQ7xsxX5Bi3m+WwyKC63yzYqri
uIXMRHyKv1/XgObE1HCjX6meFkfwi/HhpoIaifYjlCKuEdIlvCgIggfOJnAasBF9lp/61yr0cBuk
qwvPet5Lx+oAVgz+4Kb9ZvV7vyD7VgLdCjDGBsNNI5L6RSPWsng1xUamba/Kp0bu+hB2Z+xRdJRU
O2DBDYdNhMehp7UdpiG/i1/9wlmAh8lXTY7mAeq4XHLrlqSwMmLDaIBZijqhJJb0CgVR6ng6jkrF
7EfP5DQnmhCJl0TEfaZX9BzwxZ880bzwvs86fGo+6KY9qDxfH65JbEY7XUNdsSDSqkmiiBf06gze
4V+XCdYLbnuBf+hBSjwiCTNg+03/vUNXgLFJm0mKpUkUoLCOqw8n5oFWMTojMqUzgsEqFl1fCt2c
XyxLE6VsK9++pqBadSjyGOFxThpfQMak6dFWtY5rbLv0KuMMqQbEwzd00wpJxDJUI81tK7UT7ZRt
98R/PRMzbX5pPvuUVO2vS3JVDjJNrBbrWKUmJU4vbdRgFkjWaoDzgMauhMoUbPwXqmYC2x8uOgYh
DuSv70i3Fgt0tfvJ0vkljsKCvYXvKrQETzzOow1U43ZiGaxpYlTiJVqfSXnFBTazNita05XPagY/
zBF4q42QDdrgRzapHaOBNECcFwSqV+ulwZB3Dc0c+MeOtDlYfi2R9tWPTmQe0MJfJPgYWfW+6V0R
0/JcKRr656/KDzaItNi1ZzkXDbjzoB+Tf94oqPBOidHPwpfkXNArsj3XOnSdPcwcMl1UTP9Fy82M
SLq97fcE9mahgH9E/UhXqoL0p/nzAJU1AA7W/nYF8OltaH0+qDQgu4ykx0TnchBXZM/hqeT7+JFW
7+4yXU4oaTR+Q3xaYLlw35rLd3wMODjAS34LGrJsfrdYPFNIhKTsgz18LcCCiH0a5HgyTkUaYYtf
6Bb7wqg3D7onH6E+l7bCzFZ0EVIvtcaVipmCKTgqnzjJgTxZU9A+J553z+NrCKEFHN8tOWv1xsmr
r2hL9WYbBKU1mDJAF6v3EoC1EVlIPeKtm84HV1g30v9sT6WqOb6BtNBy79PlFCJO7LcI/PIWGNA2
lLugboZDFU7JZBg7fh71AhLzvqyOHYsXi+e9X6CbpQkpAYppOlhxv/AYDLCOc2etjc724r5R6fRY
SdghdCXbm2YH8o4TbLSr+G+m6LtjYPzMq04ACdOJK+koZP1fvD525WZpraP2PWBFMQob8vbF1jHj
cIMDR+RdA0KKhVi7YmdayyXXitYDFdo3pBsp6dQDyUSk8l/0wLmknXCUcvJnDORBFkboKGjE+H7e
QYb1GVTXP8zxrxzFlmayag18G9xx9DlFYdxOyS8xCGBBy8Ee7VTRnnwi3StIX+ovYbODeuFgiVig
/06+x0FMs+1GFJDlKRCxvTEm5dMzsQGkJaokFaXeuPIz9hkPXpZUxVy+4aaH1N170LBd5uMNiYPq
ZdOItZqI/Emmf9qIYdasgFpMvlJMHiT2qN7tPqGsufM4KuNZnxGgxs68dusPZd1pcpTeQPrDfi+D
5740vm/FbSmTzRacONTWnEUyNKxrRmPlkY0t4mIjC7ia/hwRaYkGyfjxmh1rTbo294YEPZUT98OG
Z3mdBeBswNri4U/ffvHSIzd0Vdq+Pev0CRrVtSmJfGuB+IHbCOGj6SLRW4clhzvcvoUMIitb1m//
yvevi1dibT+QJqM7zPsz0f79brhIh/seuC3eqr2wkhelQ5iaK8a5muaJ4BPyrUhh1RGmGoxRAteD
W78/JukVtzd1ZMCFwBTHvYK4+wjjW6UP3nVnKUDRWCfU/yJT8vFLXu58s3lteCUiE2AGTrqGKmJy
cur9i7Y6nu7LgjQNYblR5bJiWBUeqaWl+KdTfuMZkx4TWqOR0b1Yc6BSmDUru6yq4RpBSu+VGfOy
0CfXllsgpm6wVVb5PNkXQmNgUwEIt3eMKwph7P3zhdgUOnjQ/K7KRrzJKKGMJ12QzDwAE/oootAU
RgXDdinUIe11xwoMC020Zpk+INuhukGCuM86Lj2TAsRcaIbXSYDVS4QbZjM2LpVJotGicnHqEl7T
/v/DRglQRkUIYUSOuw/Gntb6TenMVfvXta3cVHNIRkY9XZ/YhuLbq0oeS6c3DzpgZwFeM6CAFXNF
/JaLPA4lIAEMA1T+5vj2Xp3qqXtJvvifj9fhaj6UmImj3v8o2mEGoaH12Pv47qDiR5i8groXhUlq
Q9/1inNJrA7QBlH9oGFqyn35I2nqoX6qK8mZto0Yhng7YzHh9+X0+8gtVzD2HB0UfOfhBZSyfxDJ
ZAU2bdcHf/ELetpCL7a15qbAfY79rnkfq8vkKbQhoLLKoUSMGA2uTmCcWHf0VltxIuEduliwOAKR
f0uxqt7IDZvqWufHOHgpx9fJ9gwr2T1QNtwUImADIZpvTwqTVts1OMiLBI0TC6lkZZfUpOtaJQSt
rStXtPXtHPlcLlJ5T2pNUB4G2U5EvqqhxDDyM5GZcVF00RCknqx0qhC5cm8EfO7xL6H0KzNvbCZT
lgLLVAtDcrIn/HyuOrlnjb5iCOeEj7JuoVtWthXENpTIU9xaoYAKkj9qqH6ALFxwGsN8Q5zf2cQC
YuDRC7wA3I30/Gd/JcxYyPOPwlNQ/jEVUHgSOXMrZ+s3Q8Dzd5EoEmBn0/uLFnT+6xEmLGkH7oc4
GpfgDfpuZraFw+ysQAY5uQ3ngDtdM2ucxbG1AaAB5n3ghMuugDkO1sBrdnxuR10twd2XJf5+BuMA
BQFVr/OUhmfON1TZXBolCi7uivw5mqBZKvItZp/p2Pt1ZZ8bCmw56/Xm29lyYtljlBXy11Ku9RG5
B/bNXwlgaK0UdkMc6TChEq3voHC2a4zj9K1scFWxVlNSmr0a9CMSinkYOztBWlGC09Dn6TcjERN7
9sN5/KjvqK3YBLLu3sdcNf8RblmoFqgiIyfReexKD2BmHoa4FZT9wC6e+fHGLtDFhS/GvEsm1dnd
MXvR1O6nnoOdo3JIA/Ff80osnqA/kVcu8pZdGzd9INwpo8NcH63OktZTdU5a25YMcNUQX4lA+Kyt
ffY/lcLdI7kvOO+33ZRIHNFwcsxTVNU2I5tP5WuQYSorcoDeu6HC3jAqFcuxPMzQF9ldPDVS5E0J
9FG4HcTaKenWf25cQQpEN2Hz9JY10G7xg0d8iaav0xx7pglZJM8QnLoficfRo8a0FcLR0wW0YB2z
yFKLADmrEtTspYyLPteW/8xXK8ohGb7Ze3h+jFrR2Egm0Xr0uSmw3I0VMsIypexsQsLGeRtJMfjJ
vBegvm1YuUaU5+vTm1+vS40cgi2RryyOA9GmBrLboawlDwbQVo9xv1eWTsNcgobLnlFU5gGNbZbN
ekUUwQBD/9VXBh5evf3Q0yUKrYdRIr9QtNbxwO315lpNktYD05cf5g/8ELeibhdcq3QuVSkAp7QE
hWBU8gNpOyffwRZIIaQiIHuOLhlVQ1SnxT4xGsTr6EPbbFz92bnhiiGFOVWni/fMvSw0BG/8UyfP
ZNNOxWMWi3qPlqTZ+Q6h1/bl28dt/7fi1Hd+p43UfB4UE8rI3LnAvBJPTF9ynpogLcaty3XE1zYl
BcUlSasPMqjvdFnX8llvxUu7LOfzznzKNB6MRV29NQ4Jfgjdc8G7GM7TKh5EFopXicFH80/F0khW
EBGcfnl/gQJXTBb7NCUAA6j13Z2mHZUJny1xQ7cQQ6lNm4whyILnMAOP5+PrYtDMt5Ap/CnhnX6t
qLUcE2/xJ/tIl2zw6C2KI8fgR0DDR5ENOMeXUH7lPLNluRftQVlgABZS8qGKiKZqWP9MSxKyMb/m
HtB2sa0ARzh44puq6tVeR2s8FjBiQmbGNX/b7ct8PVs1ImF7Kb+brbgVVBQxFKVEQ9JcAee+qzTF
iqFhBiSwuCPynJQm5+sfB9hhxcbIgxV1drWAQXWDwXvohvNSnTuPpviK786EAFvBwN/po9ExDnq4
wCzZo2DIKH+dJvT+Ld6AIZ21XYCOhx62himVktBhBaX0iArj4kHrEhrUfzRzzQLge70gBhMyCLVp
xgI6PWhXyQqtv18efvls49D39HA+XQzc8srawQ5vlAmmHuE/ELg5jWTEX/oWiOE9I+1MDUDeRrc3
JVfip+rNzuzDOnGhamobgyyLNvkymqYO/0hONPnr/2VaTAiWQqsGhdTefaxQdqagqOtLewUX12LK
C4U3VK7cZHVe7z78jkJ9md7zqoQb0BfzKklTdqV/j5G1y0wqBLqV9ZP31rdOXnPlahF+9xCnNdqS
UbyCohIKqyPRmPsnyXTZ/hR+FZGFUrlLyokq1S+ROTdUxDLQcVG1SspO6HMFOFjOtO/djfKMkIPA
7RCzj4P9Poq9ULp0eeEyO+FZIodkK1AOryKz59oD4L71Sc34yOzLrKY2JKUQ7r1nTIzUdAKLbS/w
9N5LcrKYUf6XfAigjXAomQe9IuyAHGHz/DDMgUCmy/FYP/agFWBsebQ6bjFXzALlJ6qvLHghnywZ
VeRD2+51egH8fvzG3/rzYIXCKzER7S9Z1pJdE4yV1KjNAg0CxDKmwprq0DAmR+m3fRnVS0O8nL3X
XBh6M+pFwpZdoNdcQPaiLwOM3KphKFYSkpVHojlrqIJUtYshxB5M0BrJNqmD2km6Tsn8mjGguA9b
+r9Eu5bgbbZUFIeHGm0D5VVsuy0nhZi3uK9Fimtkn5O0NRVyWsOzsqCWTq2m41RK5NG7n0x2dvaS
Su9kFf54ZnncYf1+WiIBuQ2wG0zkzTYpOhdEOHEO6wzQlE6cFTj+K8muoaOfyO6XOUG2SfWqVLu0
p5lCQ87tom5+yePdEB4vCmAYg+cbt0YOyYTAk5dWmj9Ju6zV88olNLo1SM2OBVe5EmHeZE8Vx2t4
st0W+YxJk5NFCGmXLet0YhM1XYHliUFvWGKsnnMoyA5jVYhcfKs72yZqaJNbtYQgSLrobv4N0WSg
QO56cKfGqLRaXJG3h7Y2mDftWeto7Kyap78vtj3qWwimo1PmOhehcOitKB7n7lhXFSnIOQvaZpoj
OMqL9y8d/p/7NNkSTTVieqQuNVqpfUBVUL+wJvC9Kosn5QETMLD5tkcSf8pef6VnWkIR+C2tpyHn
I8tdqm6G+ILN8Q5v188oabNRq9i9DHwCD765qhEA8I2go5oThp8lFRo1cGejYdcZWg+Ejv1tzsb9
NkcA5dNxklPVYMO44eWH4OdOkjE6SqYVjbmgLIbbpShHNAc1cvR6hETNR3+HrLvHnCrRRXBwHn/q
lLOB7F4A1z+zFP8cmFzaCfyOLrfTw902VM74MH7ACQ40schm4Gw5v47Qg3q93zRgYkjm3jOcPS5f
6JBr408eI2V8IYcpQ1YT0+8O+XJiL9qS7EY6r3lxOctNDscP7MDNCxodltjSqOmlfNBfHCZBJnF9
MEmHZW2RsVvfHUjOd+61s2Zl5UCnBOSmLENhTvOQ+HYDWqdY1fvy7E5WXkZUAJpxZ6R02zJf1Wqs
VVAjHT1RDBPgXjhUbl+iXnuKdEer9hNf6IMN+VYJad+817eE1UTZz1iSGne+rWfHCGAe9ak/vKqE
nsCFzh5OeW+ImiHALS9u5XEdGzAo6rJi8IbY7c/IArMpEnMei+vgB+uOUHnDoDCf48a9SqUbFmwx
4AjA0ZkOutkkUutgVuuKAEAKqfM/CbglYRtYxPM7R7m+eMRWzjH2m4gZbwlQGHpdXdHKqTQBWOco
5oq3Qtq/m2wNVRSLC99WeXEVx30Wd64LU0UF8+zX8kkOj6du9ar9OeJVYcmD+spJznRQJpVra8k+
tX5NWLCXanepr3brOtZDaCKU+2PqGCnT9d+0pfjUcZbVEo9VSfH05ESh3Lp2WUMYEwDic7O23E7j
3JoA7aYrECexk6FjLdl0Zny5FSYdKSYuoxt9aaGPObgQhyQdIYk0IiHX9PevouWJTuYkf0tSm6fK
/qPg5BagdZSm2C/jjPv8kyppXg7e/Zkx6/VZAfwBilE53kG3RFluke+ANbPK5BpDjT/H+FRmyqw4
vqwvpYxzMNjwrIXAkhYNWBUjH0PwuDb+W+5zb33YgIWQRqVm23ElFjsfGfr+Qo77Dcz+UCbtZiFT
NoMlofBjfsfYRpq+nhX71U1zHYYrkmG7h5S+ks8KyKW9i81ludAn3IjrHUnyzYfedjr9Xah7ChrA
I3mVLz1Dzj9nmkgqOhKUD5+PwVQ7KfbpIR3y8uCPJ6X4sxQvToTRs9QWs+Qv7uLXjyOkdSE5xvSU
YxE8lD/M9yEvsyyngtoMnkJ+cSv1OF3CoL/toHUgMb3ikW8YH/16M4DKGBMM532JadUFd5xIWuR4
ACzS6+Pk1wVquiAGlBrqAC0MPJxWRqv6ch4V3uKzYhYW5n9d4uC8I5jH9Pj6xLXjTR4R+Ne9KYI4
qY6zRhUUK2XN419xYaNbjmjWOg+a/e1FvU+Dtg3RkrNS1DI9qxAQBOCs05Hppqeg46jdhBbRaRxj
wQ53sD0stM8MP3fwa58kXTSLcIvyXAh3fsRg7qrynBK0/rAXEyD3eC4jcSVjkgR/6V7iU2LTrvf0
bcr1UGk/DQkVDBjSp4mSWKAbpqqhc8mWTld/ijNPxEW0AZO9bN/6i3jEk07BNXLU67uiXMtFYDvF
Bf/TGzrIz38kdK3yGMm9dsvRZtoq6U9WPX0mppbj06bjE+6auxvFg8qpWkO8rY8UO5d+bvzfpvgD
Q+ok3ASFt10jWKJhAxYlAk3N2Y1L28u0Y8djCGx5yFEVYf5sVW2IwiD+uLluwojRoEfHWdRWzpsb
LK9D71dX0R20CzNUu/bJCL89UFa/99HWBBnsRHMObKaJ8YGKHP75DA0I3BeQSN9NbgzZkEedZsuE
zzZqER5sY2GMlYonm8+oqlJD9+gunUgWbu7DF7OZHrhZzd3L+5wwM1oTuZHq+nluw+BPxkC0Pwqs
weqVVSr86QD6lB5iGprgc8USLfQG9soW6BwQYr6lf3SlEDAyiV8rZ0UyRRotdM4HJCsy83+A8SOr
8+F0h4YUUAfY9xMX+7wCR1DjVsQ1RVhTjaybWBN20Z5GZjKmaCJ3ckb4q/gej5E78XN2lqNWX+JP
zS5iPrzAUEqJP4NlDtEY6NFlZSc1+WCBy0EDN1ucI0mJCSppwQo4mgrfkkAfNIf2yrklQo+BYaNa
/3SnbK/1QJCqgPgrHpct3xln8ZSJ62mjjL5pLfDo4E22pepPhCl8OqvXVEtcBZS9VDhRyQ+oOLn9
AsgTwqEWfjnoYglWbH1EUqPEPgw3GYxapmX5zbgjxlCXdycEyxwzdH9u9jsyt+ACO/S7wtnAG1UW
hC9AGjhGuO1J+BCvKXxswNL0lvuL2BxsST0H5fKseQjJhWUfQQptAP1D8uv5nGIoEqhtKDBTOiGU
YsY1MLTfQCnOEDtQWiGbMTQmU0piUnO03JzjS63fkyatZQ9S96tYySHmYRtxJvSyFpgkKwz2oML1
mNnPb5rt2MJTj23ECaBI7IcB+JATHbeFKBCr3JH+NjKODj/cxUGdficg0IaF8H98Q9g6d8Fsymdg
OZFtfJ8E5cBeKyLOjSoya09GKwzsxBxfSpYnvARxD+MzfmqxaZnBKZqmS8qSpUKt4WSLwnRZEvV8
X3usNicXJE2B6Tpg0V5oYXoRcEqd+wPnUgl6D6PIvdcwR6DTHt3FvEv/4a7FJPtNJNRNTBxSQjYd
jD5wa8kGD6dY/kD9Lm/PRSJU50oI94UI4xxd3V3aG7fB+OmXY1LjLezGImEFZGllgWNaoQsIR+z/
w+Kgm8KRgJe6P9mP5Y5dreBjw17nRMrP7DtNOprkN4N3mH3jcqljGSC7xq8xG1rgzU3f3laZ62J3
uEKDxJeLKMOsnzUfKPJy+J+nRJubx+kSiEVkh4ROF8mvqoZ77XdwdCuhdYQlgAW9sSWqvixIE0bg
jej+j56XoTmkmtO6IJqm8CXTkwyC2A9PeCd9ot5MNeB933FU7jLYjWnMuuUU1fdzC7v/BQQPO+y8
fEuwUbdMhx868A4IUmvNFVtuvlm23d16+Kg2GGkJvb5YXgH15s3c4+H8GPEgcChVStm3AZ+Axy+q
UemGt7gMaJMUxY3nGG8nCQHOl0g1Tz8p4XQCsWPKsfaah5OFrjVEsMLuZwmGB/9Nv8cPxIyDnTfo
HhC9HCuZk5fiGDE70vSPgQCXHqyfAkAO9k2T268UWOkkpuydxm1fPWCAgZkzjbsjyUzz9+p+2fB0
xnMLtSQK21CSB+7cXBq5DGh6oHfCnR2U0siV8TKK7BRMOD8EQI4P/2I4IIwj33Lmz78R/lZuz4cK
aVJGnKecZroy3SIk0Nc5ivkPhEErFl6CosSRJL4DtzKT9/G5EVU7Xk9tzG3SjayiS3FA9ZmWY8+m
VaTBBDjab4sCLhBpJZqMGbC7XbpHfYxyDVGAqyOjwCbX+6UPn5OXSdghUA/rZWdm5YDFfs/t3kVh
fOP5jgfX63tKmnoNpOUcUlZcc0rua07WGU3GnHnRa0yQl6OHaZk+uHY0dRVRWxsYnte6PEnNEcxv
SJPP/+1osWUwZ34zpkvWT55/Z8fwUaLm6+BbZYHXTnMCLQvjmSdtkUT/GTbJh/BdZdf1YY/mcIRQ
IcBIb1wx9OjDrSxn6s4VHDTDwFF08MXpG7ldLQQ6CCFajtjXlqE1OePE9G5MYosZU2fRlzZy+FXT
ZFN3cdzGu5gCF/eyXDb/wLOCriAfJRKUo1FEvd9+VArQqo9S9WONLyfrqJeKuMIC8YkEO0EnBWDO
csjdlSFKtoUAo5DdVQXisiamsrAXis8DP5+yFP86we1qw1/04kZC4CYUB8/8+9h7RnF+5qMzfrsP
4NkqQIH95VlB0bYZxDk5zKO+lEuDaaul8LVOhbrNNJAnJffTL/cKsl6w1sB/LXwEqbL0R8TJPbDy
9nGVDjaxgxas31uE1V37lh+xZ4SEf9zbzVp7hbJqV7sH4R+hdbFODGOkHgabJMg0aHhqP8Ct022J
c4AWHGv5C00sXlHy9gHAko7os9MIZ3W+QImr0656M+fLbRoCexQsqz6YJQlFwkxPlSlXpBBdXWhw
PnhRUVqQoYQ8672HHEG3OKyZ1WKRpawmmSw/JLMXcIYxIsFxR1TjNuK5RtKcg2V1w87Lsq7r8MxS
w5OQ5UmtxkF9c/aqEIfPAl+rAay0l1QxbfRGvEwS38nwj7FhXXDPG5u9Mv8h1aTs8/p15VcNTBOY
7yeVOb7OUJzoh/8Z0Ye0QpGwmGsUDAZ/qQUnsgr07f9A3oSgHTWws4zcvr2OYhp7PvTfsN40qrCq
BL10NjlAQKxb0ZcxWYXmds9TFg5YdUh7sTevC9clPaGkWPq4ePa+j8rWOfXsRNRcpjzjJ139BLBu
K1E7zBJ5ZKIxBdmjTfgn00MRcdQMhfDFJnrYOS2k37JqGoxztMtxp2InwXOzBxFmskQuLy+TiwNQ
fjTo2S5FcDckvs47xvlDB9GwA4XvWX/zO2cDYStj7tOuYsMDbR3XBBMQLUd1EJ7r543bF50YUy9M
4yerSFo1ukXMr1EpilivgxfV/T4QGWIrX7WT/Nowm89EwY0PeyTULcAQoWvWb8HTFzHieXjG8jZb
cto9TUHNpTVljAj/nLx8LTa5RWzeMVJYG5I6Ww9ZU81Q4oP8SLtU2g5R39AUPL1xab61Qh1GHK3E
BYkE7nr6REkROsxyDCYOM2Rf2BZ0rXdxCAHsffB5mM1rRg0+OF8gg+DruI7PFA+qxJsinO93ULYG
gVQ+wvO+Vigxv5/slZ+Y7nA771LeGkj+o/OcuRJ+fvvOWlHAqsH2qeRAQY/n5z1maTrtYx0GE3x/
w2pd/XHFMNBUCFDZujHlzjdn2hblg8UUK0uPL/xslMvUSqIP3kfS+TMOnLmRSkgAtBFH/B+Kc2pu
TQSF2sj2xzBWd9pef7n5oh3Hge+A0B/8TCyoyDDPSeCnNro1F5PECBU2ysoPT0OppbFQyplSMAG1
K+Puiw3FS8RAIa7RuoPQP2ZOpEVSqDqbghb+Fs4B8MwWp3a4czuMtmBGq9qKrj4MaHIsQ32U8WHr
JjmYYpbdrJgedo/0Pd9bfxOUNJiDU3GHwGsw9hKRhqBR9hI//P3ldNyMH0FgGe9yhIn0DS63aCeZ
kbFp5tfmmTruqNOuSKBGm4Syuf297AK/umnOFct+H5G1baBIWcoXXzWjMMefepRrZjZWbBh4gE0Q
AaA7Svx0/sEIBkIcvWdYuRPag300hIVRRzhtOp5cJhapFCaUHbwtP0i/JB45lrWKeaGbR80Wdri1
Hul9AAXlQcqRv3BaYCBbPxhhc/fvrntuAb8sK4LjtTtM91gB/7OO8WxbGElAR+llgASRXSlyTZVZ
MrtSP2KcXvfJQT6Wg2aDxjvY+Hkeu3z42jWPREQK9Fh/Sx53dRIiwNu084ieDX6rTEtJE0TH8nSC
mzo24QUvcviMV0vBiuxD/TUWW1XiqOyKC5DxXVlENJQ/RSTomjssjcFrlDp2NhWClSQEuaUkfX4+
Q1XrJMiusFgVIW8+1u1aua51UTDq/IEV7/dztQjsJn/O2qDwgHgpQSsxb91qwzJv5w/4z6ZwJvWV
+Eo9d9aXYAne7zMVbfcjjhFv5rCzr6JnHGwpC6uVKGRoqM1QQRmXY5/ocPxfCVA7wN19ZgZDGLG8
/gr0BarP/0WZebYzUgIUKPNKY8CxE9ffNszQmlHUwEGB0ShcLCURhv8H15y/iJctKelTXU8vPkmB
ude+NBte4b46i+2PexnDMkfobu3p1GnqaIi+T7IcZFvr1rOs8hclaf245lt82ttZI6Wgj3coc2zK
kWCcRUV9hoZzVLA2nYNqpRj0X71zRhy+0U6PwhtvCeVGC9DMvJOpglLbZ+1TsbXfFfaa71TfnOKk
V1QxZwqkxQ1KUi2hSWT3J/MTwhI86tsXDDP9407LX4JxIbapA/1MXmtWAWoSqop+2BlNa9xrESvS
d/91yIk2FW9Dp5fpUCmixXra03T96TjEu+BUsHmHYT1sq6tU08GW6cLl19Sfx1LkA4PTILaC+z3m
zv7+fwU5sgQ0IZ4oRhE/2FlD1j4iIpOo6dIUlTsLtVchGEAEinuSC+ABpvhe9xGIGIIDbW9Cst2X
RTQyJ1J+ztFPWacMKlIY3rjE0o7zDuJAWSVqe3AaEB/LiDyP54A+tMbbTwLnVscHgmApsfSyknZT
LODJp7LHOo0HzbCj/GaM5MhWuOEZjUdE0yLFRy1ldT5ZqfP786A1oxFOoeJMxUnc/tJaQacpoEeh
taZO4U7Ozi+1gENjEx7Ly0+8h3QqS/P0rXa8DqKvvR+A5qye6OdWI/d46kdQXUwqWhRDwlX8ni/7
w1rAxQdfhALSlc+veQksqR9jmcaf1Zq/OT4lirw3VxmQxlEe1qytc1adUHEMC3Uqef4Bhsx7v1eD
4XgcySDYY6w1RBikAmjjOcOKPBiJb45Lxf3x3iVjK+tAe1Ffj/5dmtV5cMinWUZLtZEGIPWZ8lf+
n+7Z1X9qiZDpmXyj+sCGph7evscJlvd1uJxixhzKzFROn1U94xNq7j8a3NxbMOn1iNbSxlCYSywl
BhPL0mbGQTO1PwlWOmXApN4mrTCyC6ZZBU4307i0Gj1vUXFnPvHdL9ozMuYhZA4pCA+bKLQHZcXw
sZhLhHwoMbqpiRN+M9tQ7hFjrr8+AGExhRnuaWdcyCXs+LBd6IXLd5GwhKADR8UQanIEgXaPldpz
Fw5zEkeo0XXEO1BvD0I9xfUxjmuyvIpaj2UdJyImCPAziJIxy0uNZjfCETVr5vU6Fm5w7SX4PLH9
3ZUbpXG9vPjIA0IQRKCscYHlkQRJcleXYvsrQwd+Tzf+vvNj2sQZbOQ2KiOrMIFae86byfVKTqfi
v5JyOeNUlCFTu2rXHj+1zSXpwZv8HSQDlF2l2tSJGx1xR4Z5ceHP49XgrXmKjpD3W84UvNt61dK6
DyYb9E4srDKGe09BX/Cd4or8qR0QnWQAp8Q+orMEu+lvp7u5h/hrAT0iOGsGDVZZdvs+enc/imgY
n/HTBL/skBq0p6VOgM4c8hzHRTqNi9HVjo5NtnQfv+yTs9v2xXbAEXoOShNIthRQfHUgJIV7vm5c
lndTSI7cIC1L2ilVtcVv9aSpGoyox7SaBlFwJz3Gv0zdQqVF+Mi14wBfKfI779W1xwtTml3txx5O
pkSjGkjnb0JqI9zP0qRirKOhzKrVRNYDWdz/8qIn4SXvkXNzPfBH3FGSaE3ZEtfVk+KwAo/x/guE
gqEFwkpmBU8RNrBrE5+B3TsyqCZ3AjL/ECZgy4dCRPavIuFA0RiixrvnVZgVuHfWdE15+7XN863O
ufs2++TmIv512e4MtjjZfKGWY25vP4NLwpo4Khm36MtKxbRnL4r2vESTniRNQSF5uQb7plQV+aBR
bT6jlXoMfNi0Jj++5RFTjrysNxCf43rNWJYtJj8VaI7NZjjljIaEfCLCB9WliVS6nuTnd+986rQ6
bQ/qpR4IdcBLubsGIeMwGu7BrZQwej4GcryMQodm+AabsjWKdehPQBL6WUrwEMhyjw5G9O9BTDty
Rd4g4bz/UcO07LNNZApPCOxfdjdaJo3020yOnY/2bdSev9Y372QM5dbwTzhiA7L8OHToST2MPMXX
MHQM6SN9Ci4srx0tEIdVeOCvASvWUC6o+nUfiPjn/iXItAPwZbLRxp3zc+vUAwAAOu1N3sws6P+7
4Iq1aQ3p3VnuyS2vVbdWlMw5Lb7rp1A16T54s+lfOQjPXchCYCQIgQgydDrC8epxLZrSNqu1cXfF
3tBvU0VqFyRYgy4+k/f/tPJpzZXhZbpg1W3MHKaFmg9dyK6YhipGjKAQsPGcqzgj+C3U9x/iFs6C
6Sr8ba7NmcNlMUOuFNXmCSy/efFWxB89Y4NOHjzlxw9EErrZw8TPxMBAvkCFKwW3zhW8bDC3sq3x
2QoDeqdvdptNOGBGmwubviZWHPtFhA6aUEH59TZ4u06WDllXDc3/MZOl/ALQ5Yja/ev1xLrdzNGy
Ccpu/gRL2TObA6dOZEKtTgdfcaRe+OdNEOwvbJe02WMUGHxO8Vor2D4wRVw2p8yCe1ncFAzeQcL6
yySDaUX3Nop7X3KmNwXDty/rbF1Gzp0dg7dTeKTsWXcwkyAtNGblXeuqZaWxNLUuR64sUls96ngQ
X9kBIW8b9LL5w6aNy1hXAPZUDXxoE4LdZlds5zR8Efcq+YWllgkWUZFS6UtLxE0N+dRdPhgfZEdR
X4J99OVjurWondHqESnlcAMPCsKwEp9n31hWD6Bzbbx7dtFuDSyfVsDgJf4Z2ExcIhRSxP5GtqyA
HUKS6ZSM+A0ruazoLdu8L19ubWBnGLq4WlihJkt0RcJV6NafXL7J2/lMoLKcLIVPn4gUhczStWbQ
5RUiasJi5VyfB4hkGvPhx79BONbrdDeaCk4zrLLEtxLEltLfzCoGwBZB+wK7cwtbiWmQd28cvG25
0kq+xFF4Ub6St2L2cgOrKgraBknVfUe2j8sxGkxD5vejOBdVLreG2T3LDlPyC0cX122NgAQlJl7p
R34nsZ2AH8IITqm1Tfsmi13a0CRYCACcseXViiN/6aDSc0563zezUcXqIGUN+7K5S6Ro/5qEacl8
DM3BeFL3hkUaNxQTmchS6L2PMD7dfO5crGAxbgQFqLyW9mASsAb0nJF6HMvMV4XeO3LwaOOvP6d8
5Tja5bFO/afaReBDiKpe67JoCLccgIEW6/9jiez512K+gihfn+eOS2kPXkRaMLNxr3iaDHGQWbYw
NygG2PgXS52A7TQtaeecxIKwmTsqXKFznMvVjUJwpJ3BaCjOOwMEqKBYlMlXtbqT1gL9J3Np5Y8k
xciEd4n2MzP/T2MClzkF0bzF4dSHcZmU62DLD/2PtjzFwihbnyrIiq8xJwOODtPi02oQ1FfiAvDK
Rm6T5LzWjymbuCvOu1YkmiE8TmYnoK3XZBCdxe1gBTvumw0C7nA0d+ukzYM+HRlmcreQexk/PFt9
mtijuSITYEeevE7v2MYw4WdfjlEa4S5V53h3uznxU+l0ysMo+SdpykWbsUjdH23V5sXKrBIA5D9j
jkd4nWFA9J5mX5FXvDeTdDKSoxqP3GuQIkYGpRwqlHYBvBzs7NBCc6gh4wavouRMAVRWMc/9mqnb
9zKTkdvFRFj2Jz/I4oK3gb2vBnRzJWLacVW9h/K+3crOVcFjqWOqGV7zjouMiefUM3RNzLpRk4l1
bDMmOuPcOKFSghfaeAoK3NR75rtCFr2OPTstIwtXdT2YlX/1iPopSd+4Kv0ChabBFqXGYOY2rwy7
58zEUn3NG9CIZKUa6Ej7ENhZkBKUU0w0JfhmQ9IkOOPoSM8pDOGLFhvaUilGsxVlEYAPXzZ3Gzwp
MzsgDbgHd/lrqEOMfbr8FO0SvbZHyzGbsUSuBVKCro2QxovYDys+AnyvIRCUesEc0ju9w8LsEDE4
q06o+3IBbNOtoF7dwmArFqW3kjJ5GR3wjuM0NaoGF46+RtnO0frL70CUvG+0HsanGnszkNONfUhd
O6nYRn4W57R1bptj/CrUGDf771FTfhC8UBcQmA+sT26M8cXAyza8wtULF3DJlz1n/ovNFM00GTTL
LzfysmQT3B+moubhwOT7+eoyqstxoJMob1KpA7aoZAuhIvYJRxxu5xnSmFT5mRWLJy2amr8oxvSr
ICDlGm37TVPka2PxmoyMNyQcwKgNYRiPxVorWSlYZ/BiEnHheenm4aWLNveAzvCdXiRh1jMBwrAw
ILm7gr6ZJFk+fJTDv0tLmdQPEG+BTbsfw05j27bNe+wKyWAWWsXmFQTAtFmR0VipUGAYsYW2DSsR
GpXZtdy6uQL+nE/Lj5sFvrHcFK+OMh6jGabfIoOF2CS5+yVpzcXazMHMoKlNdXbXIvzPl8JIAxVm
hMN/n/wpQdG1l60OEtWyKSq71DaRJc7vW/rVna6uH9S/Gv7RxVsXJlzb9ZYxltydAq0OSrY5nX6M
oYdI7WmnbRv08YHSpWANVVt1fy8wNAILl24J1NXXnsoeat3624+x7w4R6sNlvVgE8eHMQVOEvXVh
cLVUJ0knYZB1GnrsQY362lxWryINh7HZEfgUMI1266VpoEZ+q7S7DM6R/9FwbXGS4AxUau7nVQom
RF5bDtk9Jetc869KGgDJsx8jINCTMg2jYeZMkuL8EY40+tc2mIvDpFSH/aLKUy8x+n7Ry28Xz/uy
Zs8yRz9Mcjt3ArGzyEsXpjGfKMr2BSReQXOS7QQ6RMLjn3VxE2rN8FdeEH+AaB1NIo7RoBxlwSIw
UEDf7A0fOK22nIaT6ac4E431lgO0lG9KWLsqTKpgTKHWqOKZFjUcXoGO5tOpgYYJ7ZJg/JJnUKSu
XOq9BmAgj6giPLHFDERY/CCNPvqIJeeeXM3BxADVKmGTZSK4wqjgO9CTFOzQv4hyZ/QR9jg+lMu4
9/wDntoIQOFphir/hqJnTrpnSWMbJKKBW2lT9gcyDAW7NmU/hVQtv7eYS68GeGLwtLTyyeSpsui+
WAZsBuPSk2sgn4a569Mo9w2qEkuIYxwiqTYEO+KhVAYqkQd30yPSuIVQdLgVYtFaqokgPb2iAX4p
hKUcKCEBKYdJkvDAP/MHPNZHJJwUDS7WiQvtJad9pRJSwXhAD0cGH2A84ugmoWJokuBE8mbtoMLO
ryBEgxmzySxV6be9t8QiXSb5N9F0P9b0YqkoIeKXXqWj7cuiKVTaDQ6G89M25iX5u7wnvJgwi5fe
S/xG1j/paLZeZd/i4Y1NC8JebKaX8IJhxHkXespEiuymuQgr7xlUarP9SGgLIPaT6b6gdPrlkBVH
hxJTWpoKS69hqu+c8MbAiaPGXZngDTZas1Xjmtiv3YeDPnPIjlNh8oGbjB63Aw0g8yGlSmpdsQw2
p4/HQtGWQI/AFHhnGKUPV80Zm0i2Ldd+dmilE3g9xKexEwoj9EZBfP4Prhvzus0iBR/ApASJ+63V
Aj5gqHFkDQf0OQ4fFPOXkzUGWzjiEhAe5p6tDg1oSBSB2n0HxbTbKdPHAzbcBoQgJyiMoQxdzIpp
Up+8RUh9210W1199THmxIAAJxFAvBFzZqAWeIMEWNUs7TkSDVz0rEDFdksUcXBwEwPv5JiPhsD9W
HYagM3jQyWw/+7f3rWN+k/U9vQl48+pZgpFX37pKmvEivVYpAfDxzaGY058IYeeAS7QsNKG1z1kX
nSZlGcutjqeyxMQjNxZOvJHGkPcwmmaLYeOsuNBEJ0sfqKFVN/VIb5Gcwj/ACrWsq53mXHtV/UKX
BiYMDQoWsfTBVMe/F7ug4hMf/lA40hJAlqIWkNxqOw5uFgFnzmlSL974LNKtdjODof9KsroZvJ5o
o+IOxXFpW2kW2VxZ6uJcUbPFzbNKiiTmjj6UBBiZ9PrX8vOi56ro3eB5hRwLNe+xnIfTYwVMIiRU
0wQn0Fk7cmiRaCHQmpQNBy+HK4kHzWCYZYNm/mKpvDDUoWFvyeCoFHu1gFA39ZxOLr30HPeXsofY
2xLX4FPYqURGY7hhWRjmmSqbKa/FJ3+llqBU/Puifoytpu/PTMpQTRXgslYCmesiuBA6BBg/zbYB
iUH3aVxJmjPftgipbaalATq4WFw43+iC7FK9bHmahc3I4ATxGJec3tzu54Q3pTU2nJu6U2J5WB5z
YPELozD1wAtSYouJmnMuDqAIW6g2Leofyb9EU5kDEyHk3qzeOIsjChuUxi5yNuOlCecxN8PEYDU0
/hHG+sIPpFkSSERoBxwFz9wTdtDIAKl48rdqyuq/uXHJkyQNLq3LrEhq+9NSJhVhCA9CuSgC2pSx
qwqvQDVnzdSYHdHwMD+4HGUCRwo9Q0Pxl1daCXP8CFqC4o9qC/6c3HFLQv9YPKeZ6BA7EJBSqNDu
2RGQTxsRCTZZNGxOScDUC+7SeKU0DwjuxbLZo6/x1lKp4/2J95SywKJYpfi9zsMtzGDSCApLgBzq
hmdtPmdTxMGkdh0KHn6vbX8d8tx7FyjpbYbX+Myjnsx/frGo1KoBwzuuGW1nPWAdnZVBBaZKe+WC
YBIYLKSUhR6tERqKi/I03+80NtfnT6lS7eBzDcG9O64dZ/oG/8ASkCF3bQ9wREELYfOXOOftGmyh
LP+k5x9OpQbywKdmDBX4wgbwzrPEmewFrwuWOOzpqvaJfD9SEvAOjRW0iGFWBttGk0PWo6FloH2D
BTIMSoKtL+xRBczdjWaSTDzy3PbiHGXsGEZ+f/crvcYQ+HiKWohjGZstpd70ESYMTCCYvrc8t+4V
5VZaMY9axVvHCbbtgPX8mA8P5h6/ILT4U8JipoTRhnJlBVSIIU1AuX58fWGcyQP2vw7UqzxkXGWY
yvpHwldCnIOTo+cam/On5jtaFpcNoH0Wz6n/ZARrtrzYAGsja0KwelF6PjNk83lWfHAeyK6ulCKm
ZWaW0zD0PXRV38GQd/NxoapIUCN7eIcXKt/cEDrnUfWU7JZQ+8VVA0YxUYaqBcKzvawgNPLsezx/
TmYEyYz2veV3u57AEy47rLkLGXgBAaFW/pwbaOuJb7ZzXF1jjSuEb5GitCF5J47upEAIsod/PFOe
h/kTBboc9Z8t1jwRkRekzAEhBf5ch68s9MoM931ZUiOIMqx1v8Andza1XLKcU5SK8oFQwwOX68h/
7IjVIdUXVf2ayHSe/tQAyemYTxTW+jKQHfmYEnQaxLRBFksEVczko99H2hmf8nJCaMWRHT52keYT
JyfDMFwm5uAbnM1tSiuWFfL8ao/Zw/nhleTERuub92kVljaDAAE/4a+zz6PBna3Hw8jpUun67c/g
RqSiTIz1RSVDkou0+H1Ui3ukfmWGqeXLl+lBhwAr8n87F8WfFGV0h8nGzqMt2sXAVbLszTm7v8qj
kDdgpGiNr0w0t5k90dpJl+9IvQYSgwe0k+R1BROZDGkAQSXKFWfx8/MsH+qp+BTx8apmP5YwTW2f
sRjuM4IiURnLM94MrXavfzvTpeIr4aMmB2kJy86ueJqxsDfwK9NSZj/dd53ZHOafCtzUSziPW+IT
Q8k2IcXf+IQdngsuPyAslOPIXR0jBrC0mY30nxocVnhWgY8But182LcsPsP/Iq3LobUyZQbq9hTC
AzwusZCFHsKePrfoLkj264q42TtyQhXexWYMiLCBCkIVNBZJEjo29kyplXuqGkdnWt2Wfr/ZB2mc
2ctIBP6yf0T6gb0QsdneFE0KIUPq+ulIgAMsqNd+P7ntG2L6W2kSHgZeQEWQTIEEbO2P2sms81oq
z7PPULtYMZh1gTzDO3rFJGB6i91YDP+W+dpXLYu9aIoXcioJqUAI8/b5xpZ3s51A/ghT2HJzq8OX
MMydDwG+DU2ag62fPUPMxDuAXDr4R0N6xm0PLKVAY6T2sfmtt8KCBMfdzI35QMKUCfsPDqYVcrq+
N938qpG60u68xxcyYHSM6wZCDLnrMmHefyBF6outHpxixK46Wi13yG2kMrCAYddBY7PmgfyPD/uN
gXVe9AOLU0xBJDGIN7I/lWIv/inRHcsUu9M4kd+MJ6DntT9Zq4hK/Znu5SC2kiwi2i02URHQynYn
AqyLmxtZrdcYZUhRmzllGXESjL4TN/5iyhV66aKBBReVuk+PYtpReOpMqGs0/dG6GjICE2YJSeWq
AwMkAhyc6n9xWqBaRakxfGOeP5bcncDJRQdG+MgZKQuySyXKlV0MBgHKNmL3GyQhsaGbGX6fu6Xe
SvMSqtqaPQ2AG2NkQFsSG/IMTrwU82PZyiBXszM6VCSy/aj3r6LFTTboTZvcgCqonij/MiEe65CR
AiNsHLnou3RQUlIQEet5eHHtgBSvhxufbfNaXYKZlnpYceD9cksd53uZhy6l/PqrzXscBm1sSdoI
VDPhhI8Lz//5GjjQVrXQLZ4s91V2hIChy7k4c7kfz+XVZlkDJMK3YLqDiaiXrZtIBdd8H5VDuw2k
2Tv4wpcffoetzlR0D5xrDLEwyjIWrcFzMFTld6xlwM1PqFK2iYwyrqKjTE+AmJ+FuVQuJVlxT1Cu
65wDcp3i956a0LgGKhOqJ74QoLSJg0Yw8jNk3wJhprJk5aAtzyryTpNSh+d3oOO/jGwzJZj6qnNA
5GPSdmtIk2mSUYWqh14r2aKK2IklCZofVipckK2EGnP7pDZBtr1k1W3YRFzXwFr4yg4PriHGyo6x
WEO5RkjGHQiuzZhWs5XtA9n/kK/uqMDDZrE1Z6pdQ1PNNklkAg4FYoY3P7lQ5+1HGfEBJ3YXPmFD
Mk5LV/DmvaFJtj9YwJHImph8rA5nqhQYt9hewsqJ4uH7wOM0CykrhT2G2Ma1byE0r/P5OEeFIoIb
fPC32T0rNki8r6rVAYengG/P7eTKn+fS9KRc1XT4J4pR0tzTwKxBcHC9/eaYFlURztHwwFZ+Meju
OMTgMUqeVW2u4FYXacxPX/UbVYL9dAxZD7BmTS7bcYJVUk7kfpYxoAGKx7cuEzVhIC4xUyIqmFLG
SAQ7bSGo24Zd+xM6XsvvVLBqv44i/JWbMNGlZ7Uj826UgTKPceWvEgfFANY//oI4py2wGDQidEsh
g3/3TudiWBI7+LFyYOVxfH49+IBGxAiv4Il3DbZDNXgcryABFOeMRY5j2e2BTI+mVMOv/LPaNkSm
+aarBMcs7eIA3IK8J5rcCjMmHTXT99+cgNqJEE4mJXedoA9ukpl1S+3NP+eAn5YtK3JP8tgjV5hM
DplPU/IPRtMBNv45XKMqAs6g3vTyH9XzSEKAyIFU4/pVJz9OY0sdnu5P6jS3hgXJLOMudQN78/3R
/bqqqxrac9uVqCOg1h1c97R5JsIbhHPlWAcCQtt5+vdymx8TaBrh4AEbq8pBk2y+QYAi++VsviTB
c1AOBpQJ8KqUMbauH+SDrNm9kOPz+nfgIRC/bgPSuSsL/SmIpG7GmYV/9cLCLvksfaErD1EUG/E0
v+Pp3V7bKg8bZCZrLJX0PZpgeZdgu06bxWSnkRmGoikLpJUuCxdz3pM+ZW4cOFnALq8ff9gU/3Ca
8nv6PiJI4IJsl7PL5p2nPp/7+i1HhTf0D4Zr8qy8J9NVeiuafd+vyFOO6YLSGGet+sq/a9MK6i3C
Q4RSAGFIRi8lKPnGmweuiQajaz1JJlGCv2KHWFrrhen6C9brCT7xXoVYz1SL9TzBLYOth/VAlA87
JGpT9qcwmYa/S7qMZH04/NELamju+q28X9cvLpddEPq4mYs9WR8hrT4kwgjfbloOU0ZiMDz6s1JO
MIU7nFdralkryWrO4ggiV8J3K8GD5HRecnCz/7isP5eny6PzlBEuOnLhZJivWUjYd2B7e5zSVivH
PCMIM6OjHdsA9iffU4mTuIWnjzaWjTbRoq4drgUEFgtkb92fKic4Gkx4c99auv+vpNkjveFZIZa6
cmp9n/qQMWp+Nd+17C9WHut7k7HfLPnDPX9RqO2YxHkoU/qoBz4wAmFehAhnANWH5qpOeYH8QaiQ
z1V5Yyn552HU9NLMTyM3GPAvXz9O2/Pittnnl3D4wlcY7lc/EEqF5poltYrkCMdFcHq4bms42bBk
7wXCf9L7ehcSewG5Xaur6JgaWHPU0+X2RIA/PcSQf8GtzSiS6n9O7JbWhLJLJA92YBsxKav8/5S5
HDODtfc+BW0V8dsnrEPge2Z5UDXr5oBDYSbBUJcTvRE3GUixKYcV80LDGOX4ry0tzKX7lks7G8Sr
R54lM6lt4OZR0fJ51vz+aXQPFDnmXS5qNoDLPeTcfupHaKJj6ppyH6etAHm3cA5f9RJWcILgeeTr
8D1E9nyknHvfCg00/3yAfhTg2h2kg3t9R0kChX5Ik90eJUbqd/boZ0XoNInFJ1cYMHBOJidcTICk
46UyMqt178xzRpg3W/LnWNKtbvjwA76h8DGrpxvz/Snu8LM0BpcMuINC5CUAg2EMQeir7EBhUmYU
DdrmtGUP/qUivuvM+aYzrwVxQiPBqJ2z6Q0PIJ6zZKCtljx/HfDTJlKFm6GLg3FhKzCFfodnf5mY
Fx8YsKynHDF/NYr+GfAzjW+4VAkoZUbZs8BYIDS7GUKHT+cjEkR3K5XofoOuHksn9cQ77pbBHaGO
qk01aUILwF3IsTJtBVkfMQ7KGGvYul83rGbsvA8wXAm0fCEccUwyaqmxmYEmyWoTiRjB8sunlobT
Tm4IF5Zx/FSMRkJBQCAaeY0d/vB7+WDNkS/kiNVayV/hdvt4baCTgZvQx5VyERddf1hMni59UIRz
0eFThdbIlGajVuGCBTSLtQ4g4wr9LTnd/CFE3HTBk1cr46zdi3FckypBP8I70d1zX2h8p+KG3k+t
3CGg+wpwE1gsjDZuyst+7MQXZwC9OeGzFaqKLpo1Td6r2EYg9Cfvbtb5azaVha5wHmHXn+LzQYcq
3gKCeFhii6J8C7lVtW/0U5dbv7dRGsL4qf05lJeFr/xR/SoHnPcoHNnKcDgCJ2W6G/B4Co06YEHi
2HRO8jWkJxxivY7cPF+ELsYZhyqUxbWP2t9S/SnPrZdIqEbwIzcClSqplJQjmvIo4PGbHPEk7Fea
ExIh0mC5LdHUfpscXH1F8qWyBkkg8l07577Uxeke1A6vNBCtntM0aHFDZe+GWkEAL2ZlLr0VlzMD
SftKuNwQ9BUhV3bakUqCZOCoDMK4GkPvd4Y82yn6KeqzCRX55YlTNxaoxCbm6pJCQtMtUllroaJC
XOXhKv3OGVMidZofasDas4KwRgdFcpA3TT6S4avt+MyvjKYNXb9XW4RhMJk3E05g5xG1VrsTwT5K
nwU813gv1DtTuaI+uVMQpqdnzO7UGlSJ1itlb/4s1B+H75zmO3MfAgd3GdgmJWFgvFL9m6AWqHUu
kmNe3BXWIUlRS7/Mwq2BVgl4FoNAZepXswJ/+q6tn2aPi5PUcHpKF26btzfSHGFvebttnN8Elgbz
mrAyKc4KbbdTWydF9wUmrwdu9Qqrnr5fzdRx3iyuqG1akT2RLFx07LjCVWMSy6/rfmnS7WvvpQOH
gG0RIHZK3Gi7NXG5qIioiMt+v+8r/mrB6TunqO7MzaTNssW8lQLeLdpv2otivbwzOphBTXW8B5Tt
jEc17K63qe6WLeL5RSMrjMF+4ty7rAF749zJq2/Bk7bVN6RfWLZnlI3MC50Sq+GrCE9nUk/j6pz2
EnbUPeU5dNIy1GzU93fpCAwMgNhY8d8zasftoTwYA0+YQOMkt+SLHwLzO9ZWoeLR4549i59FXAhV
OU3/3BQJdn8+A/MniMNKC3UAg/ssHzveFlEmez+Z4Js/UQbJUzvW9pT5EAy3bnwwcz1FFa1WD1+x
WZy/S3hfug4V2YeRAU3hxdiJZ1o7NZNKULtKHu3kbGiiEGutAExuQQRIIrHZxxjIhM9nhmMhq92v
6ut0EYysC7C+VSThksjH/SUctpMQMOMDYigioQxHuI449WL5G4sxWTFZdbx/DngvEexLc3boqEvp
e+7HEKzoROyyT3a5lw9nZyY6pyUd+R3WALRspqgu4/riJZReZI8rN0uK5JIDqcV/kYDs7mVI+bdQ
YuSKhumfHqcpvjaeFZtkpvaN1b9mPW+v96AxB6qZIsKfJUy/AUkLYBF+caxrT6/urkn+e9jxOwNp
j8g+G9vaO8FlRCTaJiFr1+GC6cGkzrT6JAMrWlIU01dZUkGhOll3NZm+83jgxo0+V7KCKVo09a2w
3iRJgQIiEWpCAkvMZoMG6bJKjvF0PC6+tNslKBq0vvr2Rut3jxi9UIEQm86AXyA70o2ojwjT+mcx
yWXGdQL0hYfPBIEsopUvb+VlByw9qDyvD5UZVG7ykBWuXfDmvRZjCO9PlOtMmIeKwbXxQqpowjDH
lZl1bDdhA44YZrRwG2kAA2KHpL/tzpzLbztrHUohsFpQdkCLQD4ahmolnJHdIXmczSnfMEXFEDY5
z47LWzZzT9toxMDHyxepfblLruYcdvNlD30sILJl39Q1d42vZXWhyg7k3C1Q7ftGbhCNTXG/GFJP
NymfZIvmorgSdfotOI6qOb3aTJn4qoIObKVkYG/8UjpejR2yrmPWAPqOOi1j8FayJW2+bf1lK8a2
qOPp0wHTZRYQFhHA4ecl9ibkrLxIF+QamsprUEAuyrkhnDsh8gbJR3dOkHx2J4gpzr4+7PGY074p
JvURfojbHci8vrMI0Oydq7mhNsm6FStU/7e4p+jEJ0A9WK8yTdC5uJgu9Dj9Y3UDqp/qWNwxfXDX
4m4WdV90lbkqxyBy7hkiaEl7G5y+tL24AJNiApRbAkEsc/R73Du72S4Yk4CbdwnUKWcjdOXqU9uE
hgrYX27lXN8StfTdREHn18ITHZUUhGq0XFc/nVE/6xU1g7+h3nimRbtKVaO6NS28RurRzTXIEcOO
HMUaHGsKHTEX7gJfuzMZOtjk/gaw+dZLxUp+b4mfBuJd2PU12LJ/m+SHddjGqMEY/4+orAHn/Ob2
g1Z/H1LazM4x0kGrOvUdrfBroPVptkOyY+ZlBtkmR/1wbjd2ojeUtmZhTTZKnhFtDsUxsvuIHiYo
nkK4gyD6ukpQdP3coJhyLJ+Y/v5ARPL7yy9IPlROn/4r3XNc5hgTTthvBkopEuhhMZKA/N9dSimS
qoqxNSsMU5fZ+8Y5RW6huKLf7k0yH1TB6bvfLNJ6MwDDhPI99fAH28jENYYqGAOvemy+zb0kmau7
cbJtabpO/4LZsSvEzmsiOVbl4X8CO8nRk50vcHPBLEGY82n+YkAJwHGfj1UdQ/lGHxeXzGDUobO4
/JGv03E1sDSc4D3mLtUNuMJDQ1FrXU+fMcrvax/9IXeFLoSPT3Y9eV2PK0ZKbohc171UQRxWd5VE
Dpi0ZPZJV/E+GqDksmUWBjfn8mjgZm+zgpbL0tBx0MjdbfP8LCvg29NWHbk2nWXxRKC8rlFvj3Hl
gnm80KMil6dm76vcFukBGt6zetFu43D3wTZh/NK0YC7ikzwxqRzq47IcuhLou96UKZE22OpCtJCd
a1+rzJt3mjOb1hdUcljz2nYcSIAN6qcNeci++MMj7MYDh3CnBiRLM6Q4/eXp5RW0l9JdpJzBsB12
K/rXobsadf2TQbG1rAsiGRDV0+imaueaTU6xcgzhlvgKiqO3npYtS/U5xQiXG3o4J5Z7MHOHRVW3
ly5jNFWZxE5AMUIAdIV+sONfMxolPX1Rh1tcy9E+7s7d6OZpko5wOkAT815rxPIq131s8oKZzrKz
LavZoby1pxByOuwLV6hmbWic9z6ToY4a5De8F2bfG4GUKHIlLtlDFkAQH0PHSs4Tu2F9c3stKsV2
zy0P3t53iw/+YV355d4lcYf37awLagbVBRW6m4DtJTwoCWidCHVFV348a6A0FEPQjbUHwVnJtxv8
JS9jlq5naKq2eRBhSuLkArluatRrUfXaQ0Thced4/2sC2lhIwAOsqtMUNrumrGiD+9f5aelnBQ5c
S2T9vKtuisNbP6bImwWEyWHIaqDKLsU/Bv+klki4yUNTtHVQATLfefEQaxWNGmK5MlHnDrTtMljP
rvsoXMVXyOJqcHDxdP9maWse+YqLzDHeksvLD3KAMShUvyWMywSomH2RInrNHjZLaLsSw8vrjACT
Z5++oGXfbD5KcuqeeE1YSe1Stdife++GWoOkUjFWQdccqVMdNzeC7cNipIv853sg5etw9FH8WWkb
ggIkVf3jdHgQfhqctu9mZ7QSZw13VRheLQ3WbsvKwCjIgVT8lPyDOtQwXXuCyTe6XL0XrtD7jwpS
PduZj+lZBuQ7V8eW5NJ/lhP7/M4Mxph6lByorvgJnLTAtpSj+U7MNtkqDHGsBwgS09/B8ncUrrCF
sK3JfVWIIfybm6iP/Qltt3JCmYEbqRTT0EWfMOS6YYsL4G7O6NUkmBdMqOF7suXTxd4TxGmkLMsl
HoifF3eqqdXRie8P3mud3eJOpgXR+Flw1ehmYUSzjLKHO+pdNb/q8XDVO/4gS9PwMg/xyblCjl6H
I4kBZ3nRkFKCkaQfwEgnF3j+uWlo38wI1ZD4gQNWOC9UZjQuXFWH6WSAYFHLvxvSbLBvKtzSMMc+
uuspOwndMBEmYQDbjto3KWzPe3419S4hbtDnsFxKtWQftANwalv5cHRWwR2bC2gX8hs5Rkd4lx+K
zTLPpN7MWeuht9e8lDfthgAwneN0GP+s2FG5O3r+cr/dGjqKxavvJ+ftQnXEhATFLN3FluQ/duOx
t9G29IgKvds1eO1xuNCtvShkXLbHDcJisx4PaDqsKaGb76SzAOv4M1CEpTz9F1hzhkrLZCre48CY
D+XXdN9kiVLxt1B6SrAsPSJPZZr2fiA+OGGdRTye7s6WlMG9nKCVvZd4xSis3ogzEXScElhVoNH+
9D8RuzqLuhiYcvj0yZUZdsO1F0bS1r8gn4amR56Guv+//+yEa4qvq6HPDE2roFcXqkc179txJQTD
Sx3joei68xQo1vmWamnSJYAM0AsAbWVrqIEJbKsQeupNeI6dprWJmYoA3R+wL+fI/N36IBrDyhWR
fP4plKKkpW0Saxe49Cdqq5qJdAdqEzUp8rss8X/QLVyfOgmqvbr2cgpR+bVTEtpGPoPw3r4XYMYA
C1ukY9Rs447KPOyFFXYSqkj1ajxkhlnVq13oitAuBTXdLzhvCnp3YTbfjf50VTZynlsbAHwqnhI9
eVNzDxgT14JWq29Id3jvNdwT2j8NU8uLLqajin4XbaLoljwaJK4meVzQp7oiMPJoep7i+eY16OFO
ElzELm9/sXaZ737YJ3eOinTnGNZL1T1cZAX+/a05O56Pjvi+UwmWqsZLsnbzDxaiD9LNt4aIxVmw
GAK293J3wUcZQgl1XTSU56DEirMJBopvmCQ2dIef5pwVUIx9hnxF9QCKXwd/Y4IizJRpr7/O08Wh
L6stltiZZgqcRFS+e8zRTrD/+TgXtn7fElmEL1szBRSFUKia9NthWTHmAoxD71xnZas6RmwFgmVp
D39JQj3U27IrQRuQ8jTuM3FeMPyUA5JZC6UBKCU32gwbksc2u2onJiT/USVPRTzLDC6k2pMMkLPk
U+YWoTy90k2UEAPgP9LbVTE9mjgpamWo7XrtgjQOmECzJ1ONm6A4r/QMYQwjSeH/FJYft+BrnHlu
5JhYhJhAp+iEdB+AP5NBZ5W38T/IgDmyeWx1fzeaDAhYLtOQulbICU3FPqZ8urk9azcZjFIcLrlS
buqs6s5Kw4xLshOAM6zMf3Ecgu5bPxk84kJU6WLoA8k7HC6rZO7oZqhKGLFjFZYT4gDOa4yh5Wp/
d1kgYxPdqU5Y9Xcbp2on96I6PZKDv1KuwJu7OBx7gMpbftikap3ABKU72SHK6had5+abWT+u/+2v
KCDEx+N5oVmZ0ddn8T6b10KC02Fa/RSKlLkee+Qw/fFBDINSKv1yCFF6zjQzQRHoO2azM5B/E62i
ecjjcywpxVSN8ThqgSHvofQihxyCl5KZ5kf+9XKq+p19x/sgdNl5HBtpxjS9mS0W4zZwscCErTAH
4kM3OoHJddlroZ/z0bipUM344d5mMTjtAbkKXO4LCUUfn1BnaVSo8JSJl8c+//hq7PIiVKeGJ+YQ
9uSn3hXo34Bp/GNA4D2WxXTbVrs9eIEO9hEo7erFI6AjG87c7Eyix7hABqZGVQygX0Tm3VCMmntY
5Y3THh98LBS1R8SHXoCRXJNHMsLfx3n/FYhikl4I1S2OjHdCy8BfYYeNCy5tQwH/YasNIVKyAyoq
PC8P6u7ukW40inZuFNNTgLBF5gf1vx34jA8SoWqBDAQh4b+oRXfMALMjfZ8RJ9SfcJRumqhhz213
0Ovg73ac79w0741XKZYmUqCOEcJikh0/5JCiHF1OHkJqu75+cypg35jTFu6Y6IvzpTtuGLNL4YhA
y/BVADh8DD6sdV/MOW9e9iwz/+25wBw68z7zeMTCAKlHhTxAGodniGbB7Fp7NrVHXm8wmwxbiYLw
iqwdUHYm+tiL5sjm470vaKaNgOY4RZgXRnei5yp8SKOFn6s/r71YfmiU4bfKfZJ2DkA/uEW+9xVk
QxILaeYX5mUHKlCgduTahZ6Wa7d/jWDrSF7UsG/0Itj7jduGx+SPMjNSHRTQMGJzWVhzmLtb6gwL
itnHDhMjn0mOvwe3wfO3wtX3ht6B0sxcKGMM6fjPKSm2hFKRes8TaO8LNGBmhnreKT+Dmf4qjIq9
t5Q9a+yco5IqOd831AGJBszolzU9joxWCcqy+02E0FCb9NEGj3GSbvtkIU1LYM5tbi+k38fxhwUA
8mJcG33R4IOF2oDT8cU318Ba8w1NkDX8o9Okxa1sqEwMOZsV608nrdXlzG/dc76+1xTXYeCDyewS
AfJkc8vu7dkDH73fe39oGgHmNYmNLzQXNF1nTVrHh61/8QDUiZOtAA3YNMftCI+hvDLm3e31mv97
1e0tgJzlVCWOcUr0WaxJeGSjft6nru709x5zg59AnASoOGMJe9BRRrWZ6L1FdBr/bz8Nssb9uEzp
ozwSAg0Ta2GA7gZeMwh/s+pRK9J4D3z2TOhx+DvqLC1U4JQlyEeXu1FZ2hDFKquKchFY6r3lMxwB
pMdj9QM8a+xPqL4wf1ckXU9hxeFXcHDeJVtjTyyMxMrrhI3DSn7kJyfu3IOK5a6z93TZpiwoNa9T
BDJNMuKvISnRXE5Y/MIkwqna2S4qDpm4HSFxxMQ4MaD067PL4Y/xf8tU3Eojs2+PQWyGkaimzjDz
/rJFBSVRdJrXMxYw4jIEjhDyExT8zacQI5UEDfI/tf+aA5zH7iPfBB1yBId1EX1ugv7qMEEMCF+n
k6Vqe/2rUrr1QTCj7ydxlV1h+WdtnlZoiGXmHQSNyWUpCyYmrI2mshNdHdnCMELfss5fg8whRRVE
naK6dYRy/pnSl4PEeeAThrjT94driE87VDuYGc699Sr/o9gxQ1ZnZ6O2IvzJYeNRHk838A5ZzvyU
ibRDpiGGzfNsZRcPgGi1zlUh8MJrtJfJ1T+kGobs1nuWRb2103aIQzqLhE1U7s1Ap4Hfh9LBwekW
3BahRewakR60BRfdDsVOtW2xi8uQy6UEj9xwBPh11b1lS2s1WXQ73+ATokbCvJtJghmjPreV6CRQ
sOK9N8XdxypIuq/CZZdIDbxdk/zaZd3ihMMAfdFqn/HBP9HXLPT1f1lh9wT4lBWPu2h8hbZc72m1
+GCBN/5YA22C2VB17k2ZZmKXVRXzyDS2grm4DBP1/bjt6JTcMai9YtHVQWH8Hoy13j7JuKupqTQw
7KYbSO+LYU6KLsAjbkyIv1IjrplJAOnL1pSoBkjkuwbkZTdg3L5n586tftKe4WG8K9yIr+SG57lQ
u2b4GGf+MnVZv+kEF25fSZys98JP4blYVsYl0UKIAGu3IK8zyZXNmPEEIVp2Hs+kzOip838W617/
nvuCrrXvKk37Bv6rtUVZOiXkB51tyCNI06vfmHt/+R3E4TL84Kavn5EefE0C1TB6oA69ohRnQ2tm
EPxaarQdgwO1iiKssTkJXORKZUmga5bm3q7d46tqHYl1MSvh/Mcccw8IP7UhtNVFrbsKj+cO9C2L
GiYefGfGP5NQS6CEGD+Ig16tgXskcwi26XCIy+9hoz54Kg7o8xerODd3EEnO1HI1N725AvRw3Czg
6qZDyum8L6kLOKQzH1ZTdCPaADyGO/etCT9JIqfAhungBaiCm1wW78sbEa/jghfP0rDZ1BOJyd+h
ALrNoztcopv4P0hBn6rgYAc2UOiBJzrFYfB/R+SL+goblXVKiZncYiVjsnM72C+lcENHiZWeQIsP
ez8SAZO8+tg4KjuxjHYjqWOyxue+3LHfuZD9MVRlFhBQtvuR/4d9n5GR9UiLBf0POnv0gSCvWAJU
KGbfsWP5D2K+qhmpYUdJ8Medhzj0vCwtuaxHEbc33d1hv9I+b+yd5tDW8ARezRXNjepBl2hZL4ur
S+fV+4BKUTKh8r8tYP6K/Dz3RgfK/JGVck9GzMKHL0yCPYSqW+QToIriwUowAJF9fIamrhxWpQCi
jZ850v1OwLKnU8aVcku4oYHvp5jUCYVd/o2vzkQ62KsZeksx8xH2ulg9ima3k+tg+wAHW1alKv28
pektAaO/NmKZhET+bMyXBGtIKUS2JtU8uTnveh2bmXVAXwRk6DJP+0iev6uZGvux+z7QWxCaTqZ/
IiwVJaP1ybS2G95GsFHXb5fDHEhG0gV3L1Dx+2hbkNM9tUIf2rF8ikMg3KKdbOoKK/h77nGKHlSB
svFGLAuSIE81tmOY9u8Bf/frim1ZfDD8EyNN4Zu2jYJkpx2q52AsENkDkmKtbHh2IQ4fZzZGtJmM
N4emnZwnyIS66AR8CgxZn5oi5UYzTq686XDcpECT3xAlTviYwwEOyUvZmXCRaUTeDG0P8jatRi7X
LRM+KxOf+X+rlOcubTw8h9HWr91o+E9bhdFUdunteZoApNLylrIUaxfuMnif5y9cFXRx76sHbwF+
7RKhELsnLDNuonE9NxZxgEAAd9z7a7xghviuzixNltAniJ+HLi/Nme0+1qKl8lQnDkulkzzLhhf4
BaylSadetnlTPhIBEF5fH4F+6GU/LEYI+cn8wpLkxkZny8yM7ZG6fepoKXSDYKl3QzaXi6ZTv0tE
ASIJXzQQaoa4D35oZpCGCKKKPcqHsnVM6GbuwZYodeIA93pqFkBoxFzw6U40z4fKD+3IPXv8aLIk
mfpjfoo0i4zH0dpnxXi1XSMy51Z22E9Uu38PwtesOBQbN8QcJbi9Mfi1VpKbPP5Zsq1STIudBMxH
kxCV65ylfVyRO02FZPWOLJsNVT8bmYuKYIrpCNKfetqqzOjYem19IHlkuuBo+0Jaq4Gj95BTMngS
bW3LOa0S8qvRxD4uqnSNzyq0Qx9/jdv2P0UwINDexRhcW38Tv3XoX5hO6S3Pexm6Kmr4jXMzHdgS
G5aNw+2eD0bJULo2My3zRh8RLItvzdy8Xq3qFNSRJw0jyV2P61hOUEFW+1Nqqs9pBzoNgRQ73N3K
dxN0FSMdChk2Q2upQHtXrrQAhebbluWQB/brGfZa2hG6ReE1XsJMWZW/wUWYtLxRvQY6ZXOKWoAt
6gKkPfQCX8gcPuJl7DfPZliynrmKhjwUDMHcivhVQmr+PZhcpW+Hm01GZZDVZAsj+UvfmBxebiFU
3zRJB7kfyp0zKPAGUtZZZovhE3aQUYW+yyr5rbvTHshu8iqsKzEqSciR+4Ve4AskBaWAmA+Q6qKN
h+pLgQ/G2ruFWod1J/47Uzwh8SaM4W+8XKUftbuBTuElZygcY9eyYtVVuhMhv0yDzujR7AuVBMqH
+/jUjbxKkDRHDap5IPVnuWeomIKzwzs7im/uI+69EcjWFWIAGRaJN1t7klPpg24krukX2W6fYyWQ
Ks24INg8gZ51lNGx/4hPgJ6qVK4VcbkP88g8a5OP6mndgBaBx12ZCsbRd0ZEoJBuTGOyGavlL6M9
lvov6FbV0bgmHhSEoDybI+FOzd/ucemRJJguDH3xeheqlmJDyqV/GtYfX9e2dAB1Fmg8QaxWcgc2
uUg5hzoVXWRj+k4AFM10FoOXpY/FyUkhtCQ1Aq3uDkejBXk7N5qlvFHfC1xuK5yt8Tqvw8viJwvB
7D/ETweCxf7CikNE+1I0bLMMrc6nW4UGIqbK80iHBfrCKKW3ZcSxYWISg6XvfFi+OrmgCpDjC49N
Vx5VA1CeiIas1uGTczxyLO2N6cNMY2/Xz/vbfmRNz7tlG3qdnpGM4vBNLWIed9Sazw3C8H4R3fYf
bMbsWjHIYntfbjhwySpYs9OWcW7vvre90FV3Z6EDqOv/I1U/OOkbvdO10XOvJTATWxy9/zXqm/zK
CMyOxLX0tA9ZDH+0zois2RHalg/+6iRKR1sTxlru8bEjld+xuP8vlsIz9Dx6qVx2VfurJZMO6sAq
axcONqyuOYl04k6YSfiubrGaZO/I+qILQXqJa9khOxl8Stq90KKIhj+xFMyEVd5BM4xmodvP0ama
AhwrX2Pn5ofUfocgpMuA770p3Ni1E1Oivw7RDZtCBpKI32/k2ZgmHxqDsNOHfutxAsCWIqn66Wit
VeCYlPIqPK3qu8AnVeCrPMKOa4H5Vi5ImQGLtznBpzbztuX+93wUnacsYMXotR4s+Ncu1GvIAfD9
SZrX9CEjAaajq5MgyPG5FBlC3cqCejnppWfs+y0HlW5p3pxeMxRFAQH/rvIgLmWNxiCBcYO+cT+d
HN+Lf0H6kPqS6aTsJCqu1wL8iaNFcm+ew/ibuavhl9uHAyyyWbSUNrbKCb7tt7P/TwhumRGDmtj6
jrjtzAZ7kbCEpi//yf+uC8LCMlnkwh3IP8UJrtvjdhbyYmZmzFKuAbgqP8dIa1Ez5ABD365EMUId
UqG/WqEjrWzT3agNpIzimu5JYHU5SH5BZTw/AD4hA/F9HNc4ykvauYy4hD0mioqqZJ8Ay2zUrgJC
kBi/fVSqZ/PluAzzMSo9sDAxsehCPCT07FHXVUHEVF5o3o0m/yK68yuDZUgGlSZkTc71KIN+suS7
shIJbt8vQSJzIllvDbxi28moStAYgp0f1rOzgwRrp/VI88iS+Tw8ogPe+/fr5zHycxddAeuptG8C
zpeA7piV3zU2Ih2v/Gv0eMRjCJBTjh5/I0uJZwPcVrWiC3BsrjD/7pSeJHSQnP9xbsB4tgzfo9MV
IThHXnrX/PmKWim5kI5f0/qi2yNfrexxzWWkIIpk3VhOylJ45gilrExhL4OtyhiRDzJuFYQnxVkY
clrG0CEufyciggtVpoLsiCOjXNj248GAN8iolm9pJtxoL5Oxhe6kJ7itiDN91SBuSe3sopaJ4okx
cAIRSYo9gvef65kfTvYL67qKMFODWokaMgAZBMuhhScgpKDd4dfRQQ1y1IY2rDRXj/0YKdL4Fa5Y
ToRenfrFXvXJ1vyJW/3zNjm4GPzc1rf5R51PvvMDwLaDt1R6of6hj6vsAUf/Ba+gUC5TIUBYWn1l
58Me6IMIYyT7rbwmrCbjohS+l/7veR/tQs6ajSR/X3CkPANQFLXEPZQ9WNzM9+II7tDzQUj58804
AhhbXgpDzzRD1wnNAJE+8HdFdV3lenvdBXb3NKYLNw36bbqo17yEfVuln9IXpyjqnY9f1fNqOSzg
sx1tuFTtwnLNpJ3+4vNeLND7ylFvQUkn76rA7kJuHArFRRVDPJUucwk2hm/e38e0g7hrl5YsEi7h
x2raR07Ou6nGclYYyzB08YcrTIryCZ1baJz5Ez+dTKc0EN85ZqbM5cfSzi+a4m+1AEbG0bZm5qOj
oXZH1dqKFEoba9Ezg84tylSaWEGe3aJwyRbmiGe3/BGpzXZTU/gGKbraJEdHIYvGk+b/spfBWcwv
A8qrgb1W0JBhSSI7syBb68qp9j3QBD6ikeyfd60uMJgW8nEQKV3PE2lZAqeeO97rXSnJ8cK5t+ga
Y6zX2C+IPcYF/37Dt7E2y53f6LYIqQOlfMK5OdUFW5wOyHW7kjZE9hkRB8JNvgkZVdhom3h/Ix/d
7WOth96aFj5JiZcIxKsBj/RLyHsF03FIePLFcZH9vrKGiOXbb7kNdEiT+S0sEPywXvyTvfhW0mdD
5aINUiqt5Nc0pnMvCpuk8wj1FWUkAv283nXUn1XC4nHGCvKxcBChv1965WDrU5HJYLkNEJWQ6OrS
QQ7DDKAmSP91ypKiqMrqRW3qkapu4u9N8CtGklSN7qqs1X/bsEq4Tg1hVroiyK5wNais6Q3CgoTR
lW3gn18DcyWbKmWCmA0s7e0txCHMUI/Vv6lIyu594ch+C5qxFA+/F5FWaonWqMb8y641u7xOU6NM
X6awXesF7G1323SEIKCKqfY08f3ge6WL6K6CF5+hhp0CKoe/y6H+XmeumFvrzfRfo/gb8KeRErAT
+u/UTbReCc1W1rtAqH+v+c2YBO8bSqvl8Citz5tF2564BxFeFum8YmTlfIu977qBaTFGrUHvDSP+
yp9Skgz1Q3zZW2gHayDY2MDCyABFYmBeZg6XRDuYiHtWFjCnjwbKZdY0gVdJt1RmEWmE8uI9tk9C
0s0aAcDbZM9gBaFcAoJKNOx1QkZePOGuLOA3IOTfR9paGdOWVIsvw3ir4RabkPAaQBZMEOswoqqa
Gsi+3KRRLl+sYxUAyZFCCHmG1AEmbtTSFWx3++QuJUcILy/88heqHW3cYW2ME77eFo/Q8GuKO8wN
cvfhAl/EtYSp8KCTbVTKBU9zImWhJqibkrJmAnUCE2bCfDuSY0Ijsm3UORIuOCfRM4KkTvTmhUno
khQ0m9t1Tp/oYYr4IQ/MIl49fiLH7CHHaf04Ht2gc+NVHRSYUlpo1gGlTppyMOW72yfDFKF+9Yyu
iHvvGzlD00i3loR+WIiOSWNldzn/t7atyyh/UgyLwgZj7rHI6gEEzurc7ZYnVepfwwRtWx49y5TF
TcEIGJ6tPtbHFTUhqvcQ/S9yI2jwTrmInWwnnu9oz3uLeiArOusTU0yBSqTxHQE0vmzGsUUCtlHf
6SXbyW0Xog9UoFXZ0OO27lejkC2Y5uDl3QOpeCy+yHgCq75dyjhWL3M38lYBpWjNayXEd6nq0GNd
CglnqpgvXM2pAijH5+AxmQ6Kdfd8K0iTsM8iEggd0kVCGQZAdLNfYYLZglXp6xNqUmKV1GXn/m6P
/ImB1WZ2Dx8yPFor6V6HMhHaeCNEzF/gpIizWPy6fj1M5bpNoguvwLWeg4scq+CD+NLG1bxX1tV8
k73WPMU3mlEuC146DuO/wxhsXIIRmP6jNDsFBM/QEdt3UNzYGctdCN/JkABmFhha/jpsZ+8ac4Sn
nKI35+rmC5KMA1wTbXyiALPyT+9Z5Dt5AJ79DhYHMZSrEc7RoK4GqqT5n3GlCBF8Uq0UMpIN51KE
IcG+h/Tv9QjO4XrcH6zvYkrgoZRsevXkY08PVAOTMC47lMU/IZKeisgNTYx5OM3kT1NTr46tDit1
e8VcdD5/oEtIk5irWyvFpgcMkcvgVF03JMh6F/ntKubfCc4b3XWPfdmFP78S/lbll8K13rLT4RwZ
CXx1hdEOwoLIL8sJ8xitBRb6adt2Fray9iHK3h8qJTWuX1hFLSNZIxWuPXPwmuXH5d9bymO6TM7D
0XmrkwoTurGlFbOwbz7KcSXWOqM7KLYNUz+7IDF1nYWUOSwBJtKof/NQZVYjuPWCaHYVgyWVX97/
An5pmJskGR30av0R2B8TmlYyd22gWbGAWo0LPC00AP+miqX1xi6qamDT7MXGIeLwXZa+YT3WwVEQ
MUdBLBeDNNrV8K3wVBvGPEeze9067yErs/m9gdPcpCKTDQy0BHUCJm9f6frQA0DxAS3/VbpyLF3z
IYLCgE3C2Q37e07HJ2ZY/s/e6zNztE0XaaD/VfAFddMR45an2ypDigP45EzowdKMSqnHe+2szjkE
qVVfuZAMDV1gOUYU3/13obns2ZRJK5rr3CsnDE4zT1jx7smki6sKPEh34Vc9RbHLghcYXdc3wWtW
4+pYbWzCh/23BFiS8zG700QNPD3ToY8uYGPF/62GOe+mY3DlApkD/i5lH01JA/3M1fkiLZA/DrQx
yxCfRAlHHQ6djP72PIbR4KwWgjvaWNOCgXW7vLigaaOcOQWj3OPlbncXe8oWoJBuM9N/qe4AeL6M
oODD60vuGH+bXv+Hnl2GF9IICsgAx6aquEKtOCElNJJWamnFEj8X+FwC3S0c/E5S2SHAk04WqACt
I799x/KsijCGSC5x4BEk+sYxX4Hkby5wlJOYJ73maPfCuHPrD/BB+i6I9/mLHqU3woLViGBOgIdm
MIYHxyU31IcU3NT+1gUClqZmKBIU5XixrqTDoaFisXqt2mLWkJ1Wiu1L3z2sMaVF2l3fka7cuQHS
J91h3GbqIDrFHHl0TxeCwrywyNI/vjtAiEMAzA9GIMxKgPicnQjR1KQjS4tj5uSygeyCVK4qKNc5
7dQ15tYA04ErFgoTeeeiLQD6kBaqjDaxn/RwEP2EeRIGs3r93vkd8EyFoodbXOUGpp7ZryBipxqR
hFREtJJH/0PaB2H/JN/FNlvZUzQo/5EVTlQh8DeyDqn0f67uvkGMuFpmdvwa+IoXryg6TCvc76vt
VJx3x50UwTTEFTA5SHi8moefuvZ2xKXGiWLmpdhlanYA4Y+Y82smnfMiUGBOGDeRC1gCPOCUaJhp
oBxeg2mze/Ym4KP9IK15iswu7GQkI+km8BQbP6ThuYu/LnPDr2gYOW2b4EwH2qC6WTDnPccUqIIo
AwkyaVBP3YjfgRda8Wo8gH5ht37jxTYr24f7dQjUpDTLWgMNCNtyOMy/HSAfzpJkWAH+RGF1tZfB
KwQUO7bZdA2jIeYdL3HFg4agyZ1m9QXu2mjQmc0RrNeeFHsxX7BnS6JmuBNaaWs105Z5p1Ki/8BZ
HI3tNgabv6FsMTfwXTDj1mX0ukXyqxswL8N+ZWEDHC8VKv9VhXzxYM0YRdq4DcoDx7jIgG9Q2lIE
qkmZo+0e6YBbwCyeyfjxhCcg2nVHsSY3/BMtuvNzk+Oi3TSOIDbc4rbqY3hLdFIQGrzD9AObwXIs
PmCZuSDDtbjbv6h3r5UqaJxMrHBL4yFVDdOB/y2lSE97dUnuRU1JacONuOheUHjiqZYaK9McIzVv
6ti2HHEWu/9YdqSF0mn7ldBYBXzpvhfRW0HvIgh5CcFz3cM+Nh/6W8ghNTCiZREznI2f/MgaV3Oj
YqQPWB6MatER9L9Ac4BCM75xc4WODicMFJCLv+EUIkZuPuhveBtoxpQYZ6vUtFP7E6HzxJIurU78
E6UwqDLwLVwCOEkjx27LhyZwY4SKQZGMbRpj65OOf6QZj0uq59J7ITkKDsd7FNAki4oVK5l5tcEs
gKj2QwLapF5TVOViYDUNRrfexddF1nYx14fN0TfWZWWR2vu9X0/tu10GzHAQE3X0OGygQHfQKS9N
wvJ/UvTaDV35Wa3h3fTMB6xrnbnmtHSVcZTdFAFosKwP97Qs2dxMsBh4j2i1uYOIePuoMa5BNVaj
ihR8C8EvBhoVORnJtwtcyd2fHO7Bmz20OaV/BME4r3+g4OnhfsMzx8vSoZWOUnEwedxMtnEVQMci
sFAr+anPVjs1YJi+Kq+lzINVImiZokLyfBUjbCP/EGluZX+4GXsGbO4yiLX19lzbH0obh6zx0gOq
gbGuY3hBCFOZDklrunM/0vs/aXqx5EWK/ttvG7ruYeJwtNWh7vuxlbVbmgJ6EpyMgvjjyzJqpf5X
OI5T6O0OCijsbBGP7Vxc73fCsXC1w1tvDcWEpc89+RRAHWj/r9PsBopuvkwyoIlXqKF2MNV5wfO5
GJvY2z8tiD9990qzxUIU3DJ3+t5GH2driBC91NdIEu46eSYmDEEtiQ5flDhN75cAh2MKRb5aCZHr
L2Nc8JWp0AEzbQF2AMogTHWXRg3Nsh313WXtSun7Ey91w1S7Pnm9f0/k2Y1zewrTqGGKLKTh+i3n
IfjtzXFLE3z/a2aGtVuDUw+45jo1PvOWUb1l5puG8KRBt0SZVw8H0nUaOniEspFw5jTbS2/pjhOq
2pCuk6yZBnqTMl0tA02QhPPXOMvILoUx29YQLSSALqU6t3yegSzDeCM30ibae4KDV4uh1IjKpV+B
tZ5F7OGerBVqAv2ipwFb1Lvbf1Yrg71xtLK8RxxTwWI6XqQe5szfxp/pqjRiklieQID3m7INZ7cl
DUK+1Sekme4FzYbFMhIdqAsbdQQm49b4TE9qi3i/+F6bptd8uLcBMj0y02+S1GAFhWMufSO05s+V
5AC19aKAllHS2Gmkm1nc7qeYbkbZx24WNVIrm6FsjxuPDoxopz5isdgZkkRU62/EnghQ+8F5/7d3
6EXSJhvLUvOpR5qRO9IvetuZJa25MSyFHEUWWlP7Uvmz4wnC7gLjKLUF5o2xm0q0WpDD0xD6w2Xb
QVAGU8mIXvElBroDLkiR2/FnuCXKfMedKHBW1WzM14g10/yCCsAgI2hGIazwnrAYGHDnrxNDPvxW
wSuwOGz3NUmuymxZdgXh5YaAg/JrI1WI9/5MiB7QZeWTMLcAdL64rTBVIu58rxVYFBo5lcy16Bkr
y+uRfOaIhfxqj0cS8lGNGbQucYJTx72p/J+iUiX4YMcuCTQezN/uu0QRX4LqXZpvlmpC3IGz+7WN
SXn5jVOQvhZAwc24C7rK8zcjdhHm9HCUjFR7dA5ptffC9Tv3QUO5IcndhfDHJf3RAas/wEyq/6Gm
WSuSkMYdwBDlPX+xJH8nbSzEYvkxbgdqu+hhB3xvXf7TKuJ3p7fvPmK7uRBmHzpGv/CtizLCJ8mm
hK8F6LEnjsvudwnsl4LH01rC4ntWNUvkRC5DmlygPdLopfGSzxED4HlmjAOwrAqt0pFk8xXFvvnV
7/otWr+Bb0a6+W7ofF7hWTWh8UKLtjuBS4foHv8Tlyzldpke9Khgzrp0wda89RSGpci2I2p0MKY1
rYVUaoIwozovo285xARQb13gM9Qp6zxA4lJytecHz7xzr3TJ5fLp7zzKfmHRFBAqe2d1V8Yp9Bx4
82GAkp6jHuwmPcYnYphKZPntG/GVIzXdUGt3KDEuQ9veee9f8oGtkNKvBpl1fvnzYwdhx+ktdBsd
vMA61TYVBPoS5TySFjDOP7jUXS+9g5ss/+yJ46jMe5CQ+H1vMaElWY8VqU7/4Jf2vUz77ThwnmAt
iJwVgUUWwDchI50Vu05KyyTbm3UuxvepwGhCHCVjBURgcN7uQ+0y+GGatfEUhtt4IDqtumPrpihO
r1CBcM23DY4LuZSK3Xza1hqxwHGpcBOFVgbKAojRNTIpjN5067wryXG5psB5fhWjTUYmgcspgR+q
cxm45V1JHKyv3PGtIe6fe1Kx7jy41Vvx0NxhMch3kOMBxg8ypymPbLxiqCFduTKMpvs0o10KYn75
anhVtXDedIQmxMZgkaujMEgBqAQUc+qckSkim5iQmQ9vKIfSptTrGRS66bftuMa+8TOj4sniOCS/
vQGb3uAr406c/0vTfcveGzG9hkJtbIOseFRgqfCcYVC6kGQfghp7+fyjVCSorcNXj88qgT2cfIwo
80zECWHPo+ns5NLG/x7qUdhBUoTpO+hmL0vV1wWtPsTV0pGs77NYqAUgveA3hxeVnw1UtaFoPQIP
/zoqp/j0zxUZ3LVTH2yQevxX0mEmud+y1hhph3iIKh+/HG7/UvciCZ/FF0n1soZGFJ1FUUNxehUI
q+vVxJi+krjjcafOeBmvvkxhbUdA93XmhEoLW9YLh/zaxFw7h6ZwstTdT5zdIM4iOFuXB6uaXqfL
RJ82+MwQQ8DPQ61LB2XIRBz6nSVJaz7fRo/ab6JUA5pYNjZdmENFwVEtMhN+A17fffUbWqkGlQNC
UbwGksaM9L4N62I7dfNaBj3FBfshJnr30O4vnogIE88UhQ8ONF8FXfLTEa57ECTrWSboMoD/xRBe
JNyDovEQgoPolHA6+hdddnneRA6Tro/Fj9h0O5wnVPn6tNW4dvKmB+Xdyl++AoDybHlfSROvvWcQ
5u6d5aiQbGZGwgAYCqVqSY/km5kvZUT+67D6WT5G8ACji4j1WUUmd23iNxAvLVNRdEjmCobCCSzB
Z5jc6Z/kjHd1dNq+Ol4e43Ssjfovr+KN1wQwU/wxx5pYM2j7LyWAB0rF3GFz2roodtWogCOaJP5+
x9aG7zokfID6FRh/m3bo/8upg1T64pBWWLVeHgzlAOyxXpnn1x1PksatPhkwnVFqqzLKA6vVu1ew
VpHsmeN9CcKJtP9/AG38qb4aui4eoUPesPOdsH/p0QOegNLnIL+aTqhWWAZVq/8dKm4YMrOA17zo
nn5gKsFlyaZ3fBgm70UHeiTYAXQdeKbemgmgUjOa5O33APs7qzc9lsgA2Bb4pUBDcHQs2eXUTJvo
fuz/VhRGj4RX92Sz33LIAjwZY9ply5oTffRRj5/ZhahE/BelM2fDiWWo67fRgdz4VgzPHdCbY/kz
/RdpixX1a7mCbgOytkpDd2HDdwuO6UhZCiUJOqL8J+MCxZvOu5aEroDClw+6lSm8a88EyWL5VnI0
HTOcYt7jJc+je76PpRo8/kK8ybAu5dTyTtJocx/LFEio7+Ni12jhImhuXKbzZx7u+vkdmqjrBjHh
Fn8xsxbkMzCYZjC3aTWJ1J9UVlI2wSkGo0SGz36rQ5cW4Um3v7dylDhYiFdW+M7kG6o1mdlbCLEy
kqCq3MtarSTdpP1BBrVNdVdMlvZxfg+r3IrgKxODRLUiHxbe3jRHXK5nn3iOjGmOsc9BuWh34Soi
epioyMJp18FjWwV3ADv3OkZyFTpwMytxJMnBT1kpO0t/dIS2YK1/5qg/q75r++KS+Me0g8/0XFGJ
bz9YTChresL3uj6KOBSLkpT0HOY+EjBrKGBdChkHvH/8fdeeo2wssvTkDs2jNJcUvTyh3YwHdX8A
FVmjwfuOG1i1mQPu8o9upEcYKoUVfNgbuImqmyzKZ8newfdxnoWx8AiZtLVU+DQU17ghFEeEcTd2
PTI3+djZsrfpe406KfyQavCUFCRY0Ax/9I2gSJU8MlPZHn9tMXnapua3TXAzmGwbWPPe0Itcgqo9
c2+vJCK3Wh4WVHiegl3FPeciKdf3VOUawKXFrwxMC8EFwnZ2HX1W1cCG0LyQF2u9DcSkhoh+xiKn
louM10qvoFN6qwg0D+HGW3e+HjZq9TJdwWP5BQPVWZkn1TgGAErOdxgo7PoIfUti5mtqrFAWGTPH
d8wAnSyzDCY3742oI3lBWQliPs5oCh0ExS824bAGBsjqQeDKdatlGGNiCnMAKQkYmV9BlI1XwnUr
IxunGmqw0Ufx9WF0qCF9yQVUCmKneluetWcYCShIJf02FMvvJnM7oHzjfpaIjGkfrrYgx/qzSk5h
s0l3S9hEP5i50Wo6rpvsL8PxVm7NmMIg1wNEE9WXqEUBncJPcEXykEyUN8PO6CddqWn5FEfeWW+M
saaZAbPNyk0S4C0jBn0nYd/Wxqg+wl2TZjX7omlD7COD+0Axz4XmFyGvmb3gGAw3tjGufKWZOUvs
CMR6ibCBaPY7DMrBvctlHW+mxUzLVlujY9+0SGviWi+dh+DdMh14stYvRqUBmk0VPRhdVv0olQYj
UES/ial8U6Toii726CCb9fOr5Zln22iXEEw9K4XHR+Tiu9NzLy/uZP1Mv/nY4vwkQXbi0TF2KNmu
LHDnOhtf0t/HYYMxexiG/+7hZk3rIp9iNGk6lGTNhpxQ+EgnfXT1APED21iHndfPR01F8HcOEMon
20QckX1vZoylBv+/gcacxbG+G1ZswcsJMQ5PQPzdTK5xhQLC8sCJGg67kLfV688WgQHv4rP8nfMP
o1+1TIdNWmaxX5ZIVdqzRuAjgLur1uWYe/daTmn6iqUK783fb8FEG8iaM1tTQ9J1BTp734iLeEDt
YN4pHd1J4Bj3LQGczG3Je6jlSipUmQdVDfHHb5nd3rU6q0Mtois7oMmfmLOa3aCpnx32AYezRHer
HTb/6LoxU3WpkW3T3olrKFxBxLxE8bjshyNDYWFsQwez2N3/O0AfHbHlnokmtHET6es2eQe9Hzwi
P+efHa+mf88Txw5OINFp6Sg8d1bEB04tKO79iPLMvMV2gMLOKJPViW+OLButmq2LdkKIrJKZUEkI
a8MusCOO8jyg6/WxyyLJCQpr8QAMG4wKKKaYz3JOJKjDqUil4n3NNzO3ulfHIT0paq+6txapQPJa
LetKgHJQ9jrtI5DQ5bPse/SqvC3YJVZc1uSz2qQCYf/EgHelrm9gQRp65ohz+lpuqb8OdfF+t1nG
dR2gpyiXY24jGE82/jo9titlSWcrKoWA7gJcABBqWbeRQ+BRrWmiWsYA8q/sjkomhQZA3K/sGOE1
8xavgeVTAYlk8z4EF6uV7JDCO9QNhlV8NU7xhf8SdCb187qTRFCcdmC20aC1iysGqBjAH2wsmOjH
WMykR4PbTSm8vh83wDsO3J3mD/mh+k0vXwZvasBLs5m8pltP6hluqqi6FbSNj2vLjRoZgdsKH1YK
NqUtMJLTKHArxpRQ1bmo8xpZR/92qCOGEb1QI+DPrTvmKYjVqVFaANVKyGnKV6BmXMhkhzlaa+Fw
wyRNj2Xms2MkRlp02u+J7EqntLAPrAWl+5UQTQWpbf2YfEyW2ch3g6jq03QVL9Xw75zuzjepaYjM
MRu4UvXXvdcYn/n2C8cY1wbhL91NgMV8JoFHg7X7SfE97/XRRk9TeRm5VIh5Z6BipZwO1K1cG8r5
Rm+sZs0DZHYTnS1lTD5mHUDTR12TrsUs33VjzS4UTAJCIDCGCk8T+iI4gT5GJzTbC5Oadw4S5CmX
jLukzlAiDewcHB8p84gBkVA+14JEZsxizjXfIwzg/PT80aCcz+0WclBhW2ACZ2JvqTAHFLVS1FCb
k/lSHtHtu6WNRolLyLbiN8+1m2IlUnFp4x4uSCgk6UzeoMu1jmpkOHBk+rLzHPDDf15KZ1TmwMBX
cGSeUUAJ2PUEILx4UOGGnpjhBHefB1CmBgwvX4dxLC9z5rJvyh0X9AsBkl+hgZSc+gP6rpaERW4M
SEPGKniSHh7R+pUdt8jLn990P3NlQsEi4traWK7KrRRdVGAVk+BO2xuqrch/qfk9e8zvVp1DdQwx
ummYBydeSLB4kEubmvkfyK3PoUOXtr3QiRsgM83Ho5Xk88q55cIgmh19n7kjRqVQd5tDTgStwyqs
RsGMwo+yEd6N2MuN6xZSNLjaXS6Pmgy8Gi/OQeymtFJePR2JTi89qcuj4PAtvNnWY7/nq/TI+m8v
OqlP8GgdCGz+BXitV12eV2U+Pm7xHtQe7T6ThdtxlxWoaOe/Y2bWQF1GJjKLGNcE6nme2UMdVj5W
MiozF6y905ob0+va5TdZFjj6Cxmbq4Iql1OtDUey/ozCoZU70vHJI7I2Pz7dmCLXidzAnlV94Sll
4YqiOH6U0xpiahHu3DIn6C480xxMWrbd6ZErwloGEko3Rof3+Jo1n1gOA9gKBIUB8ScUmSbTExO5
Z+FeQyuRbmJsrt2wOu4NYiwbHZ5RbJo74ARMaKHJRhv1CSV5fk9ujcx2kTzDTnR8AF5EjBeBA9TG
Swh/WBTJfrkmFMdAvuoQCdcFeM0WGpkoj96CYzyIgicjG5L0Z4gqonUNrGf9YY2nG98qrNjucauT
mr9qZ4rQLM/XCIfa53ZLfRV2zW73og0A6poNeB/GbjwBSDvxtcSJYDE4C5DC6j643G2YASqCsvFz
KCKRbUOVvYXTx38wOjJe0txfS21ziEl24uwNUs3e0ddXbjQ9e1gQ8j/RbPLgeVemnzTwLUvOTYIT
iKicA6MY81+MRSIVS4YPM8s9LPEqus0aidQmr8fek9mmb8gfPruT4pWnCHS3gtigLwMYw/nmW2nh
spSp20wyeIZ9NLaJg8jyJlOYBziMBjnasJsduZUs0wkTrLXvyCrZVm+1LybcUfkQGKa+pGmm4YyU
lUO5NgkZBSVCqDXYqo1boq9pjxl0Ycu5BWWiOW01g26RytHmdvj4AOQyOrBNGHUAV3wnQWBeDb2n
Lnoi9m/3Vq2LQmrT6smBCzHRu552U2klwZ2FtOoyDjRfJdPsq7llhPHNHm8BVsVtDsRH1r4N49MV
PbY48FtejUxxARvKepRjmWfKbMcWJY1UEzDbkgo/7c3BebBj7YenehwFQVftB8ZY7MHHh7In9QIb
qan/KWk5DVlFIGQF5UbPecmZLLKThZoQTyj8ort5/uOXvgYEi+t+38CTQX9+doLVDZtxdqD2a/M6
lJVY+eTlNR58eojunLBBu/igbpPob4pnMn1OlNVtjJ1zpaQ9EWM29RJ0YT5j1YiYNLkFko7jeGRh
ACzFu5iY/EQs97sDYr764gOXBA3KFYVt1STqX1YX7CTTk+Tx0uxlDpkZdWIlWT2awrXz/noanp7z
44nqK+JCABGx8k6oT/F8QuXJuHEi34T0C3FHV+2c9XErpEnBM5MTWFo9Jlz1OxhAVWBM7TBG6dfq
o4PBZR8gU8OSDF/9MWn0ACPtIsskwJzzSXnf8iDyWXXU8OL8whNrOdgMJcLDQuqCNEocZTbC7jfZ
AQ8Y69bP96PcpkxZsH9VupmcnRBIKh/T61yigkfvUYRB0Qn+smfZ1Fueb7Cup0GSlqx86cRH3sVW
/7RUTOkpeB5dHWJ8JK38V1xwzCx3VCjpVEVcy2qC+pa/pZfRQJKfORz2wFcqtqQU8Jm9/0IoWkGy
3ByQawYxQZaubn1Qqo/4mPx4RsofkXAVz0j+2awubFFQHNAi78+QQ/T8fPkFBsWBSdWiPCSKgb7O
T3BlTacA+6w+T8NEBUppPchqU5kxsLczxrNLr+BJXobIVK5hHBLchLtOYxd0LqDhD8gZ8QfLS4O7
pB5qnjljvMuVqIQ6bdPuiFhHa1EOBptI27jxlzQ3oTvGr9t2Hi/It4P+OGXGwXqUhJjhaSvPj8D8
F6llKp8gmo3JQ7fFNA1jg0FTpEmeNAr7O00sJn1Px2zJfxOCn55wWxYwUKAyo1bXzL/rCzrv9qsn
hcZo8PbDza5+gMArne9bN4q1xgHNNFvUFKFvmXNuOnTx1ey+QeOfJcP/8LsOn1O+Txp6S3qkL7Xe
uNHcuB9K/UmQd25zJusYjtcGBYwaUG8kxUOlwQa/PRsPpfhrGXWh53hgBwQ26gIBdVps/q9vGTL0
LAy8FzRZXyLr+/jKPerS4i1f78c0IAhCRd8BbEg1DdNqwb2lqTMH5+vU57vjP1jaOyKXvtQGfhpN
UJnI76pDBUvDkSSULBxoFXAQLpumzVc+d+NI87PDOQ4y08y9A3LKmysjsF30IRcg8bDy9ZSfYOk4
+ti7h92aUBb2Pf5BAwLzVQmxIe4pVh9nBrV0tz39AHBhWqhy28tec/D/lrjiCGAWKdVlAX5xkOSJ
DgE0AGXHdDgB9DIrAx1RlcaMDTTjFeQVony49Ac7AqoCZF+Kv2GKjNX31sXncanHFqSNpXIct0AL
0fEcv5sJv0kKh31jswWk+4S1l0m3VA2unFYght22N0Lzn1hRhoKemkY/NyYaRWmivIZDYAsG+bF1
0ON0Kht2Wb/P3edqYJtxNqJHOLKtlbJBmYKLpd9glIdr+usduVYBK7iQeRsHcHJTTVAZFuPiN3Y0
Xx66D771OvQKp8f3h4tK27C229PqAFHj0EVu+Le1UBoA/5xOkgUWK9eqv7nlKARbfvHaqFnUR8fe
BYulpfKxIQScWo4U5yQFTqNzASW3UGaUcKfpw/6wuGCJX8yRVVUhqTJoqN6lYaHQJlmZfn74t5Vb
t075e9LSdyfop0FvLm3QnNHl7lJMxhichAlDJQFr5VhVoTUgvtfeIzWmrigaWWRoOgxImNMY1hLk
jxNTKrXx9p7ual5DZxA8dTafjIOTq6eZG7haC5sdAubD2xPhcyhnX1UbEmdR+cgeEbegKM0Pfvk0
SMH2vRp5bl/JLzLQdvIaBjXJBRgjrzvNY25Dh/F4usuucB+jS63poKFguyN2yjRqHP0Eylq5aJVh
rj6cD2jO6uZpCpD0E4vwWjkV9KDXZFtfUoBe2NU33nw4bQpmdc29yELXB+dH7DgIKxIooSVm4li+
AMNO1WCqdHyI/saiampDPjHmN52seH0VCKxSXgtqHrY5GohYTBlwqtT98h488ZO0PvgL0rbhO7fU
aBxffWyLTAl0o1DZOqm+1CnFsFFcSzN0K9F7kbQ96xNCMxuoD8/C9Sobv2dqLQwLBstA6nZNHtBc
vdZFXMApzx+sBeX/zykCqXS8mFUh1UL/SlsEsGHbd5bbGRj5ATh7m2nRYm21wSm/kz9hH9Vh19fN
+1j5Qb+MEmcEOWbv8dnDeRWuBSm0rAWiDw/ikx6PtOTJBkObDal19afzC62qrQvJkhWwmNg75qvb
RQYlBgBC0t+4QCSZO+l3p3aXuuBYh3tWhzTiEjcFzJY9ekhheFQmkQunFDe0BpcGjYz/y2swPoWz
g7UD1euG1oX5CzlMOnP7K++OWkKLRDhSMZTx/3iSKZGcck3ViGM4UbVCmIpK3mDb7sPIsgd30qan
AJQqXl8s9yW/dVVBWRudUYF1jbORa6uDp/+myD29jn9IjisaAdNyUieO3iih1pFyvoIBmcVGKaJj
0v58fqJuQPrf6RoYViroU1vDxgUa4dOPAiGCubNZLQT1BhSrRTIcG6ELpga77hArpDfOzju7Z3r3
ABDkDrarSL0EAsFI0JBcdwGIzXae5+nSNkaxWRRjT+GJ/z4A8NyJrxjSOle37VxLrR5l45qki4wy
VQh76gZ9XFlNTTicV52ax+Y3AA648Uo22U0ln/H8fzb2NwJc5cp33aKK0/Ah6CTuKsKCqHopRunX
07TF36YRT7ACRV3bWCAPgoXRoCkVHQmsxEmrI0sXdNLnKM9B3Fm81LpiqEfsZeKpiJ40jcV6TPr+
NLLxnPU7MXlyOzH0I3InFBI8meu0nZT0vBy5DUPQU7Ch5sqJf+VhiFMGGETDL/AbywB89x5DnOUW
CubEH/Mr6Wkx7T/diKrM/MLaxx3ogitYfPVHGvYt6ZsmXdhFimLI1LN2D3FcF0kSwg3InK7sTUS5
ynVmjolzlkUHaM7S4oP92ml4uMn0CUBkG01NAp1ZMxQ1jjExXAcf7DZnWAOCPj3fFpjTOChAtLSy
TCMElyZw313mP3TancsZ3anjL66NnmhaC72eMcy1wvQJU3vk6mhwGSitSi8TYMwgGb+FbCM60Xly
FwC/IciIqI0o4VkTURicseGMM4hfcF3cJBXViyWspuLijB4zj1g9CLzkAeRwhAB718i4bkUjFJyb
0TVqlWVMHi9jWTaIUGBhV+sirfdkwfdPAwTuWHSew9eZNIfkMFC4SVDao0suQMU3KwJIS5YKl7dq
rw1QH9rOo949RaWScjLXMH9Rr8WHdowxk3RiXAAzQvJRp3FfXi1bomJ3mpFS81iNmtDBi1VGM/1b
rdKTmT/NXFbNNpsfRQkQhlmoE4Kwq95ezkH2npH8InarY6S7TlpoTrSRsj1z1UNcY86EF4r/Iysb
+Ci4OxU0f8D/aqjfuMPINFFedOoyHl5CbjaZHOfNIAZuv1YdL/FxPtJSDnEDreMwzbqGhSWPXNNv
qs4UlDM2fWQhRDFMGpg6YRKcsmMsGWm7REu58imCcaxf5IooXJDp8BkEKhBjWJpHrxHMJuEo3pOi
BU/J05huuDzalLb34J0Vd13640q2Ao1SvrXbNYemxDGEzPgxjhxRElk8FciEqi/OUuVFzT4uAHgR
ka7tLBMXhlM+Yg7hbTF59hX7K+o5qbsGfZ6cgyHz37AMEtFOzs5mjzZoHEJiZFWc+EUBJl8jYGEJ
6GBbVs0J9qMg0KRipHfYLKOq0XSssNf3zRRSElLnK3lzayr1fxTSa/6r16afEjgdLgPpq/9aLOF7
WBjjVhkkiQBteHwOU/TeETlrv31Fhka4F4oxt6OCRavxIvWR0OM+8BRIawnOgtGvebwZmwA+xH9R
o3wR0LOwJnCE24FiMfOXr+W/zeNafytkx7PUEplR+LNgxXhmBbu+0+uRQ33k9iI0RTsorTqr7x5Z
XyWpRxfEZwlG8ZvpW379v+SXtE0rPBl3JSQOMHRwFOJ1yLBx3zdp4H4KC99DqLVl52QRGe4bLzuB
Lhn9AXqjwRDE6gxT4IGTufCusiEV+quAGJ6/kXCZdewfex2QrVWk3LizZchSPfHL7bxjSM47dERL
Eih0MPFp04CEGxmBr1s1l6Fg3Enl0QTyu1vUFZwLE7PB8lTGsG4ZHMjSCweSuP3o9rYPMHCrSaw5
+JSRDy3e4KSXneo4eoxGXO19DtXjDGUn29Z7yEq4WMmKw6t3NA0D5zfrX4qQ9V528Sruf0JY9ar4
QeG5GNQf4D2TKFmBC8IWRQYZWRozD/I5LAcKn1N0aqtDvjiuPhyBf8FhxTsVG9ZkCKcGLqCikK3B
FVuD3Ui9omXPcs4LA6Z4yFO3ihsGxJ6BjCf4pythpi32/v+OtriaRs8n2OSyZJpArStzkERh0sxZ
ShXcmifXVK28plPVqLqKi+beo5jeboH4O5tmHeYynaDruRSqpdTCDK9FKT7XB/5rMHnBL9+UWAGk
JMA4+Qj6MIYdIw0sm/vMterTdvMGGOW6o7ijkb/71ICEoiT6tRysZ4gvPiDFPC7fEgvLluVFJ0iN
hY57StNoExYPR1RKEtcViI86T1TTAX7YWf8AzlGGJyCBdsfO6MkP94hi1Qx5b2tpBWlAXvPhhAmA
h49sXxhGXe/GR9bsSzkg9eifuVXEHm6cS3EM0LgSW8yLjwjGEzUcqEaw7B3e6pQf/+x1YnwFfc7E
zktJx5SXfyUaGHwRp02Ie0UYVgl+KELhV7bcv9GfFr0M3bUXwqemHxWcSKCA3CqDWubbBinhn1Q+
1ZSgUW+cDso9ceLuNFEml40BnYIlAOzPzP6Sy1800rRZ3Phxj1usX7dOfQN37Y78LmF4+j+zbxkj
vwEAqDuBuFnWgGNgK4BKfypBksiJoyrd8gUd8WrAFsVg7vF+QZO/UUHc932CrN9yWq79R3whmvxP
scxE8GzxB2l7ChT0xi9Lo+2B49U7GmIKPpS0/mlFbr1xxPgTKanw9aJ56amXxxY6iUt7Pu8rPLL0
7elzCHINb/mJj7O6g80a3BEEriM8PenN/p9xbL95Ki6qPv8KnWahpuK+d4ZRzrTrKISkquuQXEi0
F68H+Hs+DLQ7DzUT87hKkdOhwJJI6PswpBjuz3Dl/cw3abBNo8YMnI/y3oGLJlVPtBYDhrsNpf6P
HG/qtb1tB1OaMwz/ozfcA+dXK23OLMVlXuHs4TPWQE/B/3kt8hdeD/04BZlHBhdFZj4fXprkNQ3V
Hn+JSarq0YMzL/vB9YIsYemsro8ZdiBVjk6TM58lnNit79aLOD0FAsNlJxFN3AU3oWw6KtsDnZVz
AwlUw3U7GlFN72bZyuvpOyGvnmnaqh9w/1V4d6VEPLMohPUWfGPxQs66WUHIPPVBuXw8qkzZ1QEf
s/4xfKFoPGW8piFcPVrKYtVY41LKyNh86lDkNRG4nUR290lxwYnh+svSv1ZxS9lI1FjXWcpHIOD6
90l9n8TDk7PP777G/X74F5kLb6i1/McdrhAU5fpbyQUoeTI78oQcsZRZA79eBI/JTCgkunrXd2Pw
WYEXwprX+4UEsmI8sYTpX9+8Cnz+AuT5r7R9a/gKcRy5wrpym3FnNM/I1nR/V2kadXJOsdZ8ANkf
06wxhk68csIpr42F5jgDV+6Th0dSX3A5wWThYVQXr8PMvA0wBjPN00eokxPoTvltqzFss9pfwJnf
kFHrwHMpHM66oJcv/eQcRDwxtUxbT+1kXIVuKRBkukvgXb79JMn7er2AWjCfVo4obfr3g3t+MKy/
dcWftMWEjrx9yHb5xUQtFMPeEfxwywKOqPMILkg1rQqGbMKkVVuI6bPDg2f0pNwurMtVpXFpXIBi
Ir61Y00pkp8TZNs49aqdPx1W8nfjAh4bKJnznVaRqO+pNNrTOjslt9cJJ1sLcLy11crIDs0oTebo
gjX3Ynlioaoku8V2UXTal1OMdeO4jS85WgSkaa8vD/Msh4RflZEWhOrLAx/iuYZRIQhUVjnnGjRY
KWxvInkhKXrJGwNeUd+1/sGzomfNbQNOYHcbul3UTNxIGTpClzkhoRDP5v8bpxxqqtNZuLXaVNZr
DputItVN89SWJvC9/K5tawzaw1PVjNketZjJEOjNMhMQzSMlscHLpCFrZSbmSWWhoMBPHgE62oVu
khqplnh/DMRP7uX5ofFD4N+3K8BDC06k/1K5bEmMIFS0CGvt6XKtcjZZhH4/w40RW7dobGOGYUtg
jUdsk5AUoZ1bu0+h1EmMMwIFOIQIVtv9cvSDPURF2XNZictO/EA4dRmicp0ghx+JD/Ght3IxJ7Fe
biKu0kI+a9deUzJOcN5EYJR1jqUcY255ApvPndYhhYGex9BvAuxW7IdNLgWKGv/9HNWXLO2dSqkx
xzJn10rld1eDGWpjHQsXE1GjhtsfDO45+k7VG6h6LiSa21cNn+XNVRRjmTvG1KAipUJM4ro//DdX
W7p2TCFblqQQdWq6es2UDispAXuIvDiC10HKL8HPRaQpHemKs7UWcXTNybJBJ5cPUSBJDwI1rEaL
0VkWrhBDf8sq6Td6jS64/45YOtfnaXRIseOfGwqTYlfrRiWDsmAQGWGad4bK6qDNQQ4A11FKzvJG
COQ/x9zsdzNgs3FKZc98tj6QVEu9FYGlxDflvliDPIRuSkCmgzjUvUotnI5zCg7K4Yw6tFgzFuVS
VVbnY8DEyEd9GGM3R+AaipHHqPcCyoKnfj4tmmXmhN2cMRq/Z4VJasrX9ldX4oqs9m4NEWuUCLEA
7sou6chja9ye+U1u4dQaLjEv29h8Dk0LcqR0nb9cDXA2O6vOtdNuNwXzpCLiZRqXjp1Viy53wKKG
M/frlGNRqkFLzyVMDgERChqKAJYMCH6G0Y15Kza7TkkagV+bNofVO+uUKSUU56t3K1OWH3syHl+Y
N7dYDqoxuc7Znz0KzS47q9/pPXbM05ThKIP+7QnmM552GUseFYSYOiLNeugGhVSukQZ8DF72enTh
m4E/Pp9noKjf3lPXj+ugxRvKXYTkOenyFnkJvEdFMy3JRZTHowk0q9b0mFP2T42X+rI9rObhBTNq
RGenfI3SyGjPPnCLH8vZgrhjGPBiJDWK1PMZeHp7lo3NnLB7ZiYzQuIXih7HuMTXVazqGl7YxRZB
z6/gaENCJ/FFpfcbOkmGBgY0Z3+1lVom+kP5IsoKUQZ2iSGMjXO73dzUE2SxXqD105YBIN2gv7cC
HKHx1gXtJoqJdnuuyqjBVl7zPQQksWyHB3nDOnEipX5k0rpXkcgJjcz44z89Uas2MrxgIIpn/7ee
s25e8iHDE8C0Kar/J9wohZB0i1O+FCFnBHZ8YAdcigO51Q0842AjK9Toc19oZwNluSpzeU1R1mNq
mAySeYuYENpSZ2qtT7IrPbpf94t+xAprXt25DOQ/ay8ZwngMENtTF6X3UpX38sDQRvGcuU5WwAGR
OvRjKG3CVpU7D5NUnwht/mSnleCXo4QkgZ8K82esL+BQaH7yvpPZUMGzTibWYcvhjlEd2hxk8Hk7
crGiJtY7Yc6nwtKRX4WxLVnBBUYbpAkMIadkIrg3pUA3+PP2QDxEoqc2ugW4RvxeJoWtj6O2N0fk
Mxgi/oQa/GXvkSWfhNz5dNxFIv3ch/bjrjn94d4CACwfAIKdgld8uZguoBl8hZGuHte/b+w8Y3jn
OsUUpAKu8bYE67TkIUAwDBHmUu2Mx/1Go77rW7oxEPnbU3MiLko6H94lsiA2JO9chnjbP6VNbkrs
MyYPYrx8I7gG1R5z0ScuID9+fBg+Ig0a4MbxjlDTqTYWmkuB2ktWXowH2N7W1voKZCFNp8pIkF50
hQeQPt6tRv2lEXK0qzb10vU2mU1kJ06Y40Z/3fEHcrEDhFeX3AgIjV4ljC7aJZrNkKpCxfBKX7WN
+p02exXr17o1ICozytw0GjQvlV9cFkFdHxxdDfITIitVGn8H0UbdKPMCbcFwKTm/Ut1HA3FzhOTv
GX5HhndY3guIxpZKEIz7+avqgcj6k9zcMxjLq+n/VAXsvHD7q5ushdLjqTsCjZB88Qb2GyfsWSo9
DMPcoyOXrzuWqoAN7kxcsDkZ5se0th54IJvCdFVbrGb13kJdTSN4UIMmSjUxk+8zBq7hpO6sBbqi
Z68qnXOmdyKyFxCEMnX8PGxuOY/ej15S3yh0fNLM61YqUdu8NmTkYonEKpfsM6NAupoBU/EbWjg7
xH+40hdaKrjN2hWhUvGejXHyZ2aE9ybkn9mf5HBW73U25Eyf3xA6b/W3qmhgIbLef//ORHd3jKm+
dyPWcaIDF0cczY5qnSxe5yTbTei/U179eStT5HzOn8w4iMmx1ah5svXNKoLHOrZZ1ih6+bkbmP7U
IUNDLVNX9gYQ+Fcq2ndkgA2OkbDtl/A9AxHbJkLCb0jVa6kvQXE/PtrFHnE9s7u1tRp2a9iaOcFR
T4Mc8m1GChtua1M/Hgw9UEdSfLaYPmZkLo22s/dce5gqUE+F0ko2YEtoEvQuBKdmQNGyh3y72Fuc
MSDlvuXovZ5H87SjJxeKKiTw0cQYmjEf5tTGkqmuBS/P5CjSeOYEwDMq7TI+VvR8QhFy46Yr6oIs
165KqPZTgyb2X/h5xVRm6IkK9ACEhWX+/MeFDMSk7Gb2ZIG9cqAfcyQQzRI+JzuyFVsD1+UDq1li
xi6OBt9AQSMXnYjTGI1uAbF1/aS1VrU0yLCEvALweW7jk+/5a2GSdkE8k9S+R/+28dsgah5hvbeV
VswBna8/0CZvQEz9kF4VpQnESgA2N26rxqF+9f/SCpfpc+sC6gROf81b1wXbKuFSQRCPo4Y7ajkq
lYfNmEPGw/RtRSU7G0TEhBWmK/DaCeyk8PmiT4bya96ZM76iap/My5E2WvCTh7xe+SoCh64+weeE
fmiwrc4hhRb69EShYtZpT6H92lqAmlK5U/8d64S0QrxBCmSQaMxERO9UhdcFVABgHuJ0K0Vka+G7
Tfx+q2UVyW67VvrfazonUtUIrwA3QBi+sWF8QSaWlA5xeyBM1W58UGsL7183g7lbrTJ/IIvmjeSK
d11X0U3XqVJ0Jkk3wzry6D6Zbt/LLYLhwXJWO6WNgd5QHXmbMCu6AazPuTCVwlVSIqA7kkxna4Pn
oGHOjcKNA72gJS2fvcTCooufRfpL1H2EfqxOIUDXkGI2Q6F8j+XU3gMHsyTVx4cKb6zgY/tDrbmB
xRr1mdZdNk5EP2Mj2doxvYOP1VQFnQIMvIq3vCOxFmI3C9d75MLlEtE9k5HN0jDxGsfF3zoW2iVZ
bML/BTbjqtWRZ9n6Wq2pcwwUCFa0IQohyuKqtRsUL1CHJn1Uu9VgcW2Axqg9gL0ekqMkInUwYlkS
iICSD0R3W6Jr/IrB8RTXv/84fQGsgXrf6EWb12Fuv3FvgOPyQ3+OVtXeDm10PyeRfHR4bEj2T8I3
wsveGW7UX7ibDGWzJWX9rWLN3LkWZ2pMEWrBQmBcTx7PydLXYMFWaXlaGC0cpjLI2IP2ssZBu6ah
kQbrd9/RAbRBk4bokC/O6I4BajaP0q+wtgfesL/rDmzUxFLZ9dSpCa3jbp90gAudPGBuo5k+JrjD
Dr8dde/t2nJx1jc2jXL9qDuPrGZ04aE6SUON9ZPBkUG+sGjuh5k6PiRSvacejM3LSnhsZBe/awDM
WHog7qORSsIxHIxPS51F4eXfSydL8D7S5sVKR3KVhOVKM6d7avLP3MlnIYC872hqCqooDNFmfg4z
DTyq9ag7icMA2urwqDAn0nxUg0fB4qVjINykS65vKuNEs0/fVq1e3R+/fKf2rpenxZHvkuTgi6PS
0HB9Bcl/Gbkp2/5C8dhsnE95GuOfewCl1yUhcJVynMpmSfPXRYmwmv2GRD9A9WSQt/6v2KijU6nL
gq0d3G5PDHzFHTFO7n6Mal39XpQXGA42CacweVnlw2NN62Y2GgO9JDLGHuT9XHC8XLdfCMSmJfCy
McIdrrIp1ruvJVdsgkD2WuHuMtHV85ubqaAbXmu5bztz57x2GMO7/1Zn4YDbAYu/w8PsCv0OOXem
zzTRhEgyg8AkvQpnUM8znk4ZD5mKsmvadRy2jFiTTrTenLr+lahIxAku4M2F0DwqnlRG7kCq5/qm
YaX7GePN8HjpeLpofA4U8SV8eVs0YUoK07T7rQq8gWRyswHhDhjaAtR3pmI9VzUB6fZlu53cATj+
NuMuzdYg+xT2na0LeyhLBEDkVGvHDkhk+Cn9JvkxulisnLz+yjJi40ssI5Dj8GdhfkJvtmkfvk0D
VxzT5BBtM2TA2d7L1VZfmdUbCscgi12XL68s4YmE/MX2WaoPgAlPXSPgxmEyeW87v2ZRZZzbMV50
INM5+DN7N+7/Q407NIfiaBfWoMJoOamB0xl2+v1kBWXHmzx+sjoYH+/kOy6TZUndUwyuzyP+ccyV
5g/Niplo4KbQ1fONnHOaQ0Qlsp3F0hdQYCzBidZrKRs8hnxqEHHzHYDyk4O7mDH02eMZwekZVixa
i9oUrumop+OcFD+djcGnWMHNZpSG/6ARcg2fPtzExVa1BuXepV7gOa9evba4O+rteVPKqqJdCQn3
guVuDDlrxjbmoE003c3jCdbUSrNVOJP8kgL20QfljNRvg10KahIDHWrjHYaR0qgkOdkGxxwHEjSu
J3JlV1OiGcBOM341naBxehWTT6R6KxXHHr6FG26vM67taj94UObLur9ySYYTBIC9lEY97wQwfoXN
9KxHnfqBb0ezIXKtKo8owIyCHNjjWayqs8SSXb8rByeLJC+2DKCfNvWNtkFJdpuF1qR/8nw/8yLS
bzT+L/gDDgAK/amxoKahwDwyexi1WhUC033KBkAh8rp6I2CEFg0NeqA/64YTQz/drU1dnOMriHiz
YtHiV5KIiF8R32S37EVBhkXJxadom/vG6HraCVV5FX6U+4TkLUAEmSe4ONLjC3sQGuC/+NGXbTQi
aRJbUT5u5Zvfn6f76HusKlfcfGKOkbeFLUdPCrKJzW1Dn0JfekvCWPBzxdt922g5D/nMtsOjIDV2
K+NtRrZA3N9y0S2fCCVCWz2k+g3jvPRhp83IsvZKwFbpUmllCP00htQk1eREppVn+amdB9ghSzOI
lySrcNRrdnCIZpCKgulE5HAs6Tv+Cn1NIaGcnBrifPtJSstJ5gnd/04qccm0lOMfb5gv7No6dyZR
EEHA6PJ062DWHFwtoykT0j6DjW4oK7C9ObHjQdwkG9yX3npqI0GU4HU9EMKzJrkzOTI/5xK46fQm
WFLm6bmXefugvf+86MkT/VNAj//dsZz1rwm5CMExwao7AcshPCq0WoDAiv3B/9/wIs81nWF/faMa
TQkHZJIgihkTnTbRQZ3F6fSPlxxQlqgbLwzSn6bI4z8FLxczD8sGXSdsCXW2uFq5D27+xck6YAEg
6yA/eBvekDnEGH68gAdRfG6G/yWgtt7rEXzL3ENnpfVGQYKTQwPTdiYr5pVMsyJsw4LLn6y2dQOm
kiQFANcabxmKLOmeZQ6L6gYCTzl8miAjn/6oc2/i0aNZuNEtp4/+nEM4DuQ4DlmUpoxgQZTSLdE+
YOrpyBxUUnuOd36Id6YYbApPGDTiD1R3KsBVd4pgYv3ydw0cU56s3jMINk9FAIBjJgKxseNkx/AN
us3g0vJ5w4u1GXIFNSHuB+HbFh8v0YvjsVc1d6oZZgLUt4H3/6Cx0TGeLwiLwv4ZAWGalBDbe7o1
f17tptOpO10aPVwxu5vulgd272IGVOmuaxQannmNbb2+Hvj65I4AKotDN4QARi347mNGPNGOuyIe
7fM6JF+wxZ1dQCZIPo1+jrz87WBYb18ermI8gpaE5ktHC0KTDsAico0AzeyzbfP6a24+0rhGUR9G
K/0n+1/1tQuOX2QKuN4GoXJGC3YbeXuBwNO13pCCykG/+bgrBfxMR82tz1zjkaNcKtKj1AX1X2Fo
zc5AYeGmqPhHs0MrfZU+mLtP8QiJCjnHwx5KKdOQIZe5vxlhBn8gj0SEm90rWpyMt+BbjRaqpp+J
wjr55Xn6AUCvqL/F2udcMtzCNCZqC5SgzqjLRmbv2V9eXSadij2x0VEmMR1hexhgrABHvwAghj7T
7IOg1OGBGqY7WDnT+5V2jJyzh8aN6bnCyzckSQxnYmF66N8gikwIkURtZL2Yudzb9HsajOrMzXHN
i99mhb9YdCm2jbtZ8+neQ8bEDZ+4bhZCF4QDVdu1SN9/IGLm5NA3H6YQ0LSDp7CnhZvxzP3ALKul
g3zFYUmaewYnWI0QgY+IrPH6w+chHvbQ7MNMHWad1/WQ8sdtORrB4C3j4P+YDsG3ap/Agvn4iv94
9f/VmF6rLkGNfpkFnQ6xaFDjX5LvEPaARmHd24RfFCUBSoeKJN1DTA243x2hamOFALvXvnNcHKD5
YMwkmyhGIHcH1aT0tA6+K0iAzc7PEqSnSdy7BXfjDtN0o34APhs0YGR/RueyghO4deOWKu8OGzMD
nGRs8xlOdy9C6+Fg3UtMLHKQzYZ4Fpi425Nvj93qoGS1CII3CtZlIqBqzHKEZ8mNw7vLHejPqjrk
6updkp6Xdc0ZmxZJfAteg+5QlG6yLL0ehpP+OaE7zdk1muvQUG9IJyFu/KZ07VLVrdPjBGYC2aGr
OfFkd7mvVs6kSEnirt53BoMS0uTTg6NLR8isxp7oPgLhQ1Gkox1fam9/+n+37LnjRgUre+MOOB4t
k0OkxWSnsyyqsTKEytJM+X4CkDto5A2GWkOfRMbfMcVZjkuME+0px9m+B9ZM3C9VwR/488Vm3rxr
5l+mIF2vwujJbJ1sFMIEH7D1vlfgDYbgXCG109giSxo3Ktebo6oidFmunaGII8x/C4qcN2xojWTO
NSYduStI+O9yIyJqwEBhV+RikpQBwrDkmat/duxohpbSK3PAQU2MaoNi1L9DsQoZznyHkUwsrGBp
j9dJRArb2QhNmSECY63dLsf07V95nj+ZCfkrVLDxo6E/e3nJ2nFHnQMXfM69ZdPaAOW5nB36yTeR
iIaG9shDI7xFonQMLrjDc2i0W6rqyLzGEj4HcUcSU7fHQhx3+mvJQ8r6DoiBuk+Jqokjf/BgWHgC
1MCPLIJb8/E8haZuzv1u0hVkMBUL6bdJ/vAdH8/1msLWPWe6LBbK7InE1k201bok4StVkNDH3w2E
J0vy5xfqga4ZP3UD2LyyMKJkAXGK8Q3sg7f//s1QzsHKBPQzTpp3OaDITz68FkPUqnNnQqrI62Sq
simHrzaHlOQS6l+gAMo+2xHim4nUr2j6xlOvZHWgVZ1alS8+Xomhm4YFSfaZGdo2FAG5Nrq3JV1n
QtzKoZY6cLqra+Bel8jeLzrEVLsKXX0acnBmRKtIR9SR6YS1W90e/UNsR5DivOA3nWpKUrPBph+Q
beXnMD8qslbqm0bQMZc8400XPn9jtJuLXreDKTBXSR8X1ivHGMp2ZYWRjEbctvAxb238cekzdKj6
og1fgDWxGchsxUtifJFBMNellIzwfX8TqoKB9YEp8ehdSFANyoWMnNxt/WLoXmGIU8GdRfMkjUhB
cxEBPdaBnnuhMFOVgzFaLNTr0F5EompVdfLs7S7yPPHRUOkJcvKBcMDafUn6uOgZ0jairxVB44Dw
zpqZgZr44yo29Qn8iUTNqAlWeMcst5cab0xx/7+aVnggz1cXVhjnrVu1GgbmwrNVQCpbfRx+V0vr
uLTpaQgx05hSFY+567/dx4c5LdzQm6GHVzhsG6iFxhpF6a36Sd/T/SLNWaFmiMN4W8YyF36ZtUwf
nFTB2ym2EJ1i/f3AniV4NL3aAsJe5xhHLUOLM6XBKFnpBKn9q7WcwvZcm+9uyue6GQswRCh/kObL
FtGNxx9SxekUbGARaO5WmF+B97zIJPHMgfxCVPfaNVAdws6Nk05fiHyI5FBxhl8o8CzD6KVimKt7
e/3MImXvdBlqWhgt/lFDmKgtmxzoc0t2LF42qvDuVmddbUoNJjAl2wevzU1GYnFacBp2ViBWArhN
6lrfANUeckA/NF1ncxg3Db7/bAkylcwIgc36gXRIYdBqT0InizmfXTXlbq+Jh1GhZ1nWCuKdT5lO
Pq4wg1YeGrnTFBlyD+dDlfFPQ7B1zws2DkJFKo8jcXOx2OaIa143gDFmN3w9TACiqM+3hpOIsHGq
B1Zn+9UyoLkLOq+2QZfnOfYgS818tGWegwyMwSJCy1Fk+03+5fG1Ddvchs7aCq5p5FXmSopSn1yb
iiLv+exYjhxC3xosDn4N8j9Wc/IWcW1arYfXG6XrVjIFPi1gOh6BxyDGBTrzkJpGjd2P4R/QQR+s
io5FeA5FKJ2ocP3kMiKoXCnJ6l0u0owjeCak6/WQFMrFe+/bZQKLd7MmCpQ2yreyJWplqkwWi7A5
PA8uMCb2O876IkPnZYm/6S62RNltJO3D2QyiU5xgMc9ZbKEKAI3QHPkf0kYK/misSw83J581OPhl
1M4nXQ8aLRGaiteZy7c0k+HvWH9O1hqZBMxlOw4guCuqgvoryILnCot1or77+PISk0Lad/9+ZNM0
WZ1TObfxdRR/YlxXYwoHcncWtoDt9JfOCj63kvMOmbuVKXAq5wwQC7CGnzOvmCAUdF7k+nv620iL
EWe3RAVPaBeWIJqUkMsugfoVKNuJ7a80NnRKDBVa8xQRJpFlD2JwLhfiMfpkDk3dDkpccXAhYLLZ
5usMu7Y9kVUMADviRwpq99tQmYSOFUvDa8tQPGj44JxLCMy3694MuKiaJNtAnliyPFaFybbA7LRu
ViM66eOexHYT/4iQkjGSC1rsLhI3jCEDWGyn02MAqAL7dtoFiITQGZrhmyoCPvVV1DVhyv9DS8Rp
0ulL7zrWmvc8TrK0v1YIWyffZr9ZuF2HHG92iuCCfrld58xd4W50Wdm5/YwjBbgYoCAIyH+OZ8bS
DE4DA221zT1QteCFxfTj7SuuS/aMYKtAmRQMiSjx7X8n2k3cvymhgEJUQ42AbZLDquUkxJW5ecI7
8yhY5boMahOgvi8YLJWFk2XX577497+9AIYGQ8FwaleGxpUlqerXEzEgrvKcmYzdg45sozoxVU1r
9tFqaB10aGemCKpoaT7YEwqYzERJ3AjCrkMDKtMAyRW5u/1bqQ6l4D6fMKmcJByPeWfZBUpU/0cS
+GNug8B9rvZKTjNqMw6OblJ4ZXqbW3U9t+7NLVvrWI4GBfra3zu2T/l3prcVRZ/Eu55UZOOcBpht
HsYAYKDgYFtHcbzqLQkVPx4TSMA0x7fCGYuDq/k6HOWJCiafVx0SM+cNDQ6lhQd4VGP4imtDhL0w
HIPLmUoOvTWH44AFxM5528xToS6oOoEPJm82KL9zhh/IUi68FajNAiUnm5d8fsd6E33y8xaKswAY
GLJ6PcOUDQMEOGi9q1Vt/CGmyrOFdJ9rKALBWrHYh6rnD5IMtMQ0QBK7K9KTKKOLMET76Svg9B6/
g4zrWqTZDPKsRBvGdx7uzs/f0eRGz1RGM0mVUJDjxWN6iPRqa1Yff6Ii8iDKu72qFVAvzC8BpS7W
/MMLLQjTi2kQBNYJ045x/WpZXXrS332Rp3GlTFNi16L8EO1yvPqYvTNPNPNffi5qOt0pW8pcFMuj
alGoC4h7Jnzpvnx1CqG/J1SZt+CA8LieFo+Ku8+XPVGWDHRQV5sUXGjAnBlg63zO5gIzwSzRcx7z
qKsJq3gSAd2fJv2wCCIqGcxrVgfYTQJrQD+ZQhHn5N0MGvr+v+ky21OhCsFne8nN5lKKnY5DJywD
rZAl1+GP8tK7n3SZyqfK9fp8lKQlGYcAnPyicibmxphbEbZ0FxsetR5uojNE4AQpFPyHE2bSpuuj
6eQ3IR/MJzrjI0vDKLb60J86wS1+YGOKOoSSMiwslcIHwxFdcEeuxc358t4VsNXsNyG8RSdM+lEw
7Hvq94ccTCA2Diex3/eNZomkm/zbxTRhHnbYK10zYsHEvfaKE788xrOIMr+/Ie9OnzEd4zeolXEA
gUhl5/vOrnZGgl+BNy93LTidReXNHYapwsrSHpmGE4sxhCxRUEfH0iq+0wIDCqgMnExbsnKQ5+J6
fR4IB8vyHJl51dkYB7CIat5/rYG3GASNtMydaPLWtOC+VjCt1dBjAsCWkKPBjjI95vAL4o+wB4FA
hSuaQwmDECABrBjW04hTFEAc1BoDXYJgrXcrfCHMVtrpuyDjXeoV28Le8t2OVM4VUVu+hgre5ifI
/dwbJgxQqn8kb6/PAQq6slBAl3Z1GvTotbQtS3HkyhZ4B1M5cx/pWT7khmsZdqRCLDISpnaq1h4h
xVVXjp6xvWKmiDdRjqL2WvMISx3Al2esTgwtoEg4qQiv6EZ8hd6EKDPUuuuaHGcO414GZ2YV28wQ
SZIUNguCivasdMeRu1kbaQciaKDLjWyNgchbJy3xui7IVVtBY5X8AOVmpF3IA0FLiTFf4JOaHHR7
2++/v/LFPPWvrEgTH28GGc33BYmbsnGYiNq6SibdBraDjjUT2ziNyJ9H7VH6P39RId8MYmCke2/W
TDeOfmgf3QWKAaA3FSYHGeb2uYXJ1og4dZmxFFvGnlICfegAwIKtnWgPvVAT2RjftA4bcHKtxA1w
NNd5pI55zEZe+a+ZvAnPlN28OoM181sVljmgDap75uU/NHvD9j/Ls12X0ICGu9z4mc83I2OR3B05
c6tv0mD3YIsxIlbZ7xPNoKMCBU1NabvfufPReY129KRI0bjoIiAeS/R0s2k+7pjTnMywKtVLL9M0
miH3ZLg8buumJ8PBz79SUhmlkpFombPgsC8Eyumwd6pkLHv0XLQQAOizBYqx8de/caLgb36eFDi1
YNyqb7KmGhNcLbPfDG/Mciwk+mMY+N7Tj/i53M7acpAC0hP+Y7w45+pqyE9Sz6W/w4wSezSX7fbq
QlokYzX2Hd3hW0JYRWfp+JxxC95+ROHGo1QpQuSQ82exHCt/moLRjjvdw4x8BhyABgPJDw9Kdu7b
YTJYQa+FN9McSROPK90hfQsFC+5eX+w3HWLpgpcenVn5wdmKokAurR4Eh4yj2J8pzNbZ2o/10yjB
6UizzjzGC6ckEIPfUIzrHbO6lq4COErM5gi5vpJcxhE2P6FRNUZFbumYOqTu5qz6uWgWWYUdESwB
5Kh9H56JjekJH1s0dSqJADTn5U0fpit7dKy1NafzK4Jhrv9ybYby8gBS7ytx7zVg0MXsIQYw2UeM
ZFtIHD4gtN5m1m2Rp/zO8iU3nWhI5UPrvT+R1XTwg5gpLYLQ23ZhCVwJBo1lrwfgm+Gn7Cwdc0w6
7hJa4GWBTs82ffrWkWfPpCrZUiI2yWgsCHy+QhkNozn6PHeldjlMIIHz6jansnSHIOOmU/nmv/LS
C6ov8YJzhbBy6QU1ltDBybpQ1OzwysNrFUtZqBzi/D97MHjbPVSLMV1JiOpdWOXieqvUOK4/c1XN
JysA0xV3955fhO/MBlnQ43cRpEm+Yf0n5eJvVGCDE3kk6xJzhJHdFA3Agl/ijjSzLrwkDCrq9UzS
2eTlJ/iFe7I/J6ukKLrXtJmdpm2Bmszhs9bpcQbvSj5Hg79BOelaee/rk3zgr2SO9nttJiAL4p5K
IHAl2IGmLBaTjn7z+Ta1d4ly9xS7ROWXbxMuYTpWPAWoiJ8qVedxDHCW+KdidA+jkjI3G2VQCYrV
x3XdipKJ8gdhj29tBAS8Rydl0CXIGgMJUiY79byygzwsQyjdUyYrSO9jc53Bla2nJ6yTZAK0sU6J
2SowsVOMJ5BVr4Wml1BQDSnPPFYXHvYKL3NcXRFh99WdLK6eG+n8vfCKwXDleDXssnBdIW2g8KEq
CKj8BLUA6ehx8Qr09sLnU1QNBfR3RxenQNxT0WbEojC912qtDrVva0x2uXlrugwCb39iAm4zkZld
rLxQr1KDbXHSvUgDey0TjZze3WLKlWmzpGAt34+wNyExBcGuOsDI+nJ1b02yVXahhyL6pt6lg+YT
zU7YTUsPEsmdlR8J50jOb9aCxHo4argp5P5mmmo/8Io74yGCrJrQvpEB190IzsDRbFh1ye+fH6do
Q4MPGYqLm9cHBtEE/fy5IZ/Xp7Mdz+iPYewz82YEpWBAnuxesCFPb22TV5zvAZrapvLDtac3MleE
WPkxcNouPTSqzxBGum2iY3LILxF8GA/SmAjuQeN3yCiwOTqH5eC2vmCdX06pcZzPfzJfbNoYnlTH
Wc7Q/uNAOWI6+In/mxLSY9HaaCNBMrPZNN10UCbfcTK/KEJzGgw6jhiW1RJWtpErzxwEH2ksw0nC
baZyXgAtRETkylf/i98Lctj7bHSvRQr0Rv73glQOEzNorkc0GvUbbk3nifolsjVX/X8qrIJaAI3x
cE/D1QTf1gZs2ycGgcq+p+Fqcv5F6hk2ThQRAfChFQPR7DQZualvYTmMVeNmZQ9IHXWqBdZVLU8i
+V83ScmSk1EFL11dIESx0ei5avUugdSQbDx8eyu2Fgvgz2UVmxOUhsoH0ykg4Pp56UNKtGThEm+C
2WpW7bYyAgPgoW8pQHQ/jK6LKppneneiB6pYCzsowbFAIXhPEDGjtxMnyYmM02Rk7af1RCyfhCt3
iTIR/U6fF4EWkdDzckJezBGJ+hPPu0iPipWwF/ScD1Nb2qq4wSev1K+b+YtswIHUcot1y7BQcHDT
xk6RHMbxJPjbnPMYQ1hy30gsCFlfn37IgzEb0BZj+hP2SotknW47silrjYSsqb1eIj3SssOeigOa
lVOkl48ZuYwoffY7zFJDd3uS4i7odu7QDHq71BT8vVawLqLMwFDJljavTxBIkNuwFrhyqtYvokjc
0VrLFVfgLXJ7RcRt+JKhjWpO2VtFicD0wFETijC/gGIjVVXw+8K0mIT63Ekm/FcqdDPpVOttXwJO
s8fnNMe4zhsLtUMI5J2b7VukhOLC389JnYbnq1jrRVnaqQblHLRmx3Fm/KwNDYiOYH5wDDsebYGg
93KrNF0eR0hssHmnglURggKFJEoEcLKRu0hcDifzYJj52ECrlUJ1k74eThONsUnJPrpPzFJkV2gz
n2cBZRu96s2yUIEUXihDWSra2GtqCubWADwKXKscqCMTFBcd7fbVwTvu+KLHUQMwzJQpwWiMw56Z
5PcblBUsZflVOgSwYTkBcTzSoL+MsWUG8cCEr1LogXSr+kxGFgEcVkMIfbbJBeuXGonyMzDXZVMp
1MwlAspyI5KEuTK9Kq39zAWFqZ0MuIilDIxCzzS+uF+xavr41QushIJXROvZnR2JVJzcdGAl7GLV
aZJyq3u8zbOqd0AIbwR/ODftUNgwGs17sZS8TshIau3WR2CuV8/oV9pcW764pwK1yD9GyKlXQnph
35BXO4k3DsxQf8LGR9axPFdiGhRp4M8zuD3GYxjgrjz+y+qmzTg3lq8QCVVkmb0vlNhOYTkBcJEy
W63OwEvJRE+ekYaT8ZpEItHrUEmpDHcSUU/oHDES6s9oIr9zksk26VP8+3odhnnkmQstWDIxJGxT
wt0tSgZDfcVyMouEag1vvQfEaA5XwejVnBZD5HDhAvQrak4G0CBbJ1i77LVGIFr7nsBnnZ7wJaqF
oBZG3EeRFrjXdLV9dd6uxJWwJqfDJHWhRhcbcBHsC2rM4r8zlyjPxyWvCXYE/zLo9U8miiSzJzkH
uzG4NCwPDWtgUj7kbm106WY19ktuvRpoURo/30h4fLqNybfHfQyVP+5eVidWF9JLJ9PSQubQytKm
2sT9gqEZBuhaTQ8LwYb4KkgDlpCs9xBDtiCK8w+U5F1GN7xbu6NpfURw++ifWBlMfAIm+3/whGZv
NjKaHao5USSRUoBKCEe4+q36weXq8E2HKBDDCvfUmhqKWpXoqmyhfHV/6ZlDZEUdKOlMHAoQ6m63
0WPfeDo6bJElDWK1Xy8KV5S4F2CWkHs0DH3G5nsww1JM9n/P/nfJIz+sro0co1/K2x0RPVFxbmWX
12dQWGo37AvQE2ocN6PNr5zBUvDxED47rtzxQKsPc8M2VwM2LYbfzYr5+0nyPiUeFdFfe5VxV9Oz
qQ/2qTk3r/GE0hBEd7feuwQxoLO7sucDtQnLdzlCjaTqEbrOsdgBRy+gLQg4QDh827nUq9o0CPMy
lGreElB5oxNF/Yil3WM45zJxzitCiSuoDvaOpsVbzOERKr0nAtazf6HzA5kC9vrP93MCHevpcHTh
Pujd5LG5UCHU2fuwDmARpZZCNwTkJ+vL518MLXXFcTiBo3m5lOn6tdg3UjYt0rGmvNmdhzglhNH+
BT20GHHfl0JBzcYs2JSgy8vYRatMtSNNcNo+AdQZkb93Z6tb/LcydmU8B4bO740NTPRJTrkUk9T7
xMJ8YC7S1FUrVG5pzeM6o8rjmhrDVPIT3UxzWA2yfVqipOQpcZikjq3frL7qOvmvIZ/mNZBZU1q8
UBD5iKPG10DeOKPPBe4f1W37DkFfBo5jtFnFgfJNO2ETKwJ4CxPwvuYdL+ShSlOhhOoCdgXTQmZJ
8Kij8KIVcSPWmO5nNIE4oIx2bYsQbYVmctDuvKtg5O0XaSZeBb7wVsXak0Y2sPwXBGJpLVZdx+8R
PNBLLx9W+O2ZJrbXyQykx9OGW9SnD9+ObSr+RcL7OFIgnJi2hsaQld6DBfM/mouhiMWOejeDHpxo
wMRCtGeyynTEQrPmdx7KwYQoXua160ihMj4U3oaw5ArZhlGoWAVX/z7HyVW0nnPeBj8OZ/v8WHnx
nw69snpW8shP8J8v2aTJxn6UahV0Kv6FnhEv0J8uzgaybTNXYvhbkbdDXzzcYmhXB7VV9sJzp+mg
o7sr/nTZYKzgjhApDqPDxu8ASJCFSdx/rMHO0CEy71NLiDB1LpM2G8YbUnwVlXdmTEIBS91xXxTa
0YJ+yJ9xRUCFrPF/iYlS0CvwEP2uLpKOZCQjiPoxS0lHFWM4roIdyi0rTAhqxLr8BU05kI81tW54
5DslzSv6jvdAzeRfaO2nzwHU/GCRJ+9VePrmTeq2Atd7RMasyXvwsYI2Rawzrkia9OvKkW5vgNJj
0TZ6U/drCSra4UIJOKvl9cDFgNCDQj9MforI3X+PoaZ06KInqUnzss30WN6AeCcY/igTba+9Dz8Z
kQgUDxoh6Px3dsuYl1UUuTGByBgSpK2xmY8qHpvO2ETDv8QusU9/hUZ+N9R4zAruZ3XD6vi75BTI
JYx5pJ+OBe+3uTjcBgZ6bABt21DlFkTOq0PEEhi1P2cH9rwepkEmBbmJPskbhEFX9IGHnInMSpfh
NeIfOsv/IG+nb4AeyrtYmEo24HOefpVQIg6y/05Wa6bna9OCUAGQx2QcZMz/Ckn1WMrssKR2+oTi
iqkhk1RgWLxcW9a185IbBaqX4lCwRqW0ytxTcOlMcf9rIIO5SA8Jov/ufi7YUSFvDQHXCKQ97Ad0
zFInu5tGjDWWiboYM2k3kE7XBvUJ+ff1CvN6NTAplliFX3118N+5cccoKVOYcK1F2azBYdWhEphs
VxUuTLX7nOk6wvHEhNf6IDZGNlGSpsJyqa5Vk5Nt87/28lfeatw5lEQm+LETeRt++CyUVvWZKEch
HB6UQwaEs7bvpx1GXhaglAFFsWazGcRxk2WhxXE4Ml2C1Cd2a7qRPzEnTPPBP47jh5irSMCAUm94
9LL4Xbzdi/5ujGUFsOxS4kZ/VjHLJj9ASnegnkZ2s3XPotaN9DHRE0izmAIM5YgjePQiiNeFhsTN
AadmU4x5gadI0UN/s1SEH5MjQUk21ouIw7T11dWIWC621mJ0DzxxeGNs2+xLG//UcdF2HRBYw959
Rvdjoxz96ZkFs/x909m/ZtzE+/swCEZFKbDjuLrGGcNtx9pp3/JIepKvPj18wYROc9Aun0f3xSIL
x8fSp6ZzFsxcJjjzTB6sR5jL61W8qJCJ84V6PTS+O+fy/vJ7Wdnmpqx/6ig5mN0/Dqu7AsCPHPSS
D5Nh8RatpurvbKordyT5SBUqcMF8qn+fH+0bsa/US7Kj65qGD0hyOcVi3OjEBfQosMCywh25LuDC
7tDGuLBGwiK9eP8btMI6w9MqnbyFWbZ2g5inirNTPoUoKMneT+OI77Kd9NXHdr+XlTw1oKIyNSAa
JCEMq+oXKoVsUlPc7f8eFnZ88oT1CGmb6YniVbUXgkVXxJKA9mhi/llmAefRAZGWvpy5PdX4aa1n
L3ssWIRyKxkjkBzTrPU/oOSSzP8ASjcuSw8RXwDoJwd5kuJ9l1Tj9FMp/49f5HumWdkpV0rfeEiu
G5SKw9mbHxBhGEshy080wyoipvPLU3wlsVJZMqPP2sid1leFDAIL/cr+RC68ue/4EO2PV222scIR
Ha4i5A2XnabiL9IXoNCyX0tpalpr3R927sbEHtR+3B1r1Vf6SIdfNrnjPC/lWUYqlq34L72NStB0
3cceM6RR2mf46xgXxv6wyoywu4G1xfWaui7dn5UxlSCyApqZw/rxRQPMbpAvs0HANj0b3VorV7YD
ryJe4TLcCett1h68rmq9KTn4zKLuTMS6zVNlYGpuhA8K8kBzXF/pccEcEZdevN/+r9y6WCiRdtzb
/iKn4cogsVVLJxQ4WBiOvetFKI/9oa1/MUfdqCkZGJ6q3XSV3N5vjb1Jh/EYnna6u0lFRvCU5TrR
Fha25GPM2EH+4BUQRSaaiv8aob/uA4Wv3vhhz4hVHBXtwdjYfg4+MvkvK7iErIKQFM18QVFL5DmQ
nbu649gvJ5sS+YW39bHcZ37fhukmrTdC9E+cj087f/2RL8HDourA/2lr9onYCohfqrhZJ5+Cvj/l
rzQ6WCDApN8H4Ww6ihv9E75SrJxlqcVnXQQEpzZpu+ELYEhYNeYBRaZhnP56Yt73xIpg+fsJlSAD
GSmc+OdlPcKN8HWzz0SGnSD1ACKS8rMQWRXJ07qtcBo1EsNxCzJetP4dIjvweMs1Q83LvzLAS/fr
rLnrEEHw1/rL1vrLaqmSFlyvzdbuOz0HK07tflP2A+FIFi8VFyctFD3ENBSQwc85tkZei0PedkPk
yikn2TSRvWwBQwBskAUH2KUM08wLXCSOdayHlOEhGWCjYSKvyM4TYTVXuzmi91vpYqamD7q3yTzj
T4W4m4G52nSzxmm+PI1FyK/fEN1Q6AjRSJaXBhMev7yxE454KqEgWJWg+9JLv/GxCcIS68i+Qnj9
cosp8x7w+f0s8bdoDq8JFyyEGIWZ2HEM1EQAWzNSNgBySFwzXaXfIBLpeSi3J8O7+tD1GdBHcSN+
y/CfKwBspWKLd7alf9ApNgWLYArS011addpMP9exXqERDnuF2O6x6ewcIXESMgJs+j7XU2h6BhMx
b3C+I1cwjnvC/aCuyCmBpA78YxUxLr4PjwPc3w1qKZeZ7FNqDUN5F+s9egXXH9eft4Ft8Dd0jz86
Sym81Hh32dzIktQiFzvZsgLmD6Yqq32ZjOzchf36WULgCg55MN4IfJKZfwQhcaDehnyb5IPn4Qck
vmSjrWvUL4QZa3bUzT+20hVugkuF/gCqZOjKRyqL5yd1CwRkuMY65VIauKvpBXo/1GB3LsbDlV3Y
qHZWEwXKPipDgSOlEUHlyUU12Kix+FRNDQlHWwAMabsMVyg3L+eBYp+inYt2pJjpbXTVYuGK4dsq
G9y7O1iJaRrxsefz1DKflc9aDPHdL2J/UXm3HTceVJyu6MbhE8MCxydrqhQwxrd3XZhHCU+c2/EM
mZmVyMRCY14dorfvpWjNXPIO1q76aqEq9/IUdWK7JlHHTDA4SiLMl5kmzIaaQGGyrRPnGN33vLT0
jJ5Uz+lGS2tvo5YrRo0OS4Q3nquoCDIon8be05lkeF0BCOfUDmLIa90Pw8G3Hafmo9hifc2D70Ni
TS+N6PSGU7+/VlKDGnPkUw5RLOARx1JVaSLtuVoJWsf9JOyaEeAer0prMa773oM+WT4KXzOAXyh9
BgfH4wwxtMA7J66rr5dlUEzc9hKFCMijCWu808OaT4wJr5fO7rklC2wvTF6lKkou1FMOsBKOc/UB
aYjDlheruN2FpQGDbGsLSch/Ia/g2MCUmMLw+uuy6alLS5wlc/VexB0SsRW/KE0/IVHWd7txU5yu
CZgjzBVyAD6bVd2viPLq7CdsJBFxCd0prKrUXhx4KVlXLercbMKAJJDpRx89SY0SfLKJTOtQ3u8y
BQ1k+5cGi076zL/QCjk1RmH/l6mHZQyCj/ngM1n+DEOCiD97blMXeZMDnf8qU87b6coivAQZKZ2h
lLG0JsSKYAx/L5ZB2fyk4KQZiKFDpb9/kxHondAPvLPU4rlMjZHeRyx0ibvxvdMV52Q4OW0S2Jxe
EVhYbACR69xJsGTLvUpOHEksYtQt58RiOUsxrSZtlxzaHflYJVrbh3Mkgkpos/DFFS44iYX9uZEs
gf1uV25K7DmpIIocj791QLO8iTVEhsHTKqBnh3xi3LjhasmNmr03wcA0XLOtqiRmcFvlj10gSBCX
9NFkX3gcYAuNhw/agTk4vZvjMVG4qtjshz3+yrH/836rCp15oYFFBefGOV+0UdnQIBoTsD4y7BZP
EGoi8TAS14sVJDS3VIKP3WRcHnrh68SU0pGGfdSR9Sd9K4oorkrqt3TQsEcgaYBHLFHuGnLUkD/v
7BTbRPLPkanHDQZ6m6sbpKj9nfEP3TmTZeRWG2aiqY9VObpMOB5aPviT1eCNGQ4sFFgquejfNf6Z
l+DYbjlFzEKfMTQtES8G6MA0PL6czMfTOCPRVyuT6U5k5M30VY/hNEV9GMSslpN4MM9Sh573pqHH
Rx+Pg+h2K1dJso5HAyQZif5nzABxljlZGiIyvwtEkLJsBLoFiZnrRL0yk21WZlh4/1ZGy2ym+iDQ
ofQOcINVXlClEaI0xRut/DgxbzqQpOgKvoxyyjMxitQMtaB1iKsQIKvtrmbtW5sQdPqPkst9d6Ux
BC809Tae8lzqIX9VNynNulNd9Ur5KG32X0kqGpNsCqaU21PCxZX6q/NrbrGdvUFz4p3hOhc2DscH
rgzT626UFY7WQjUAg2Vvw1qwIKud10I3+4UUmOQVSmrXbzv2qKPsSSu4Pmp7R+3q0by8LPW+u7tG
JDkwxUTXiE9/io6ZCQxspa4jI/NopHR2fcxAheCHFg6xfyquQQQuED7zU8rKhHG0sVC+8YqcPKrY
8qhJxzhRQVLHRueFSRPp/lL65EO/LoeL54XMZjpD79AgVUzDilo4BDuzHRjRneqvsagE5Sh3RFko
GKun/pykoaWEvPsAIci/MJQzmBQ0gtuoIPSV+tVYlIbQuu9GYOstpCFefTDF3M8b/D0va3334K5i
3j3CVpQy3V81b6+lLscUpn7x6praxkh9x+ho9jT+NTSwYnCgIpULzjayfhKB0EEMp3akWNIdusMI
BrLH4zdgdALz0ry444T8Esbqq30iDGQ5dvTIdEujNStTAP7Bvqth9SvgHR41afZB1QRPGt9feFMe
lNdxWA/czIo3C5bMWkTvfKbuLVHs5ZiqLSjyWFgwW6/fH5dZneWSj0/xMaQ2fmdcCCpg4O13rtx+
TfvctUvNbOCq70Do0ljNMAt03R6GMNDfH6K/HduhaXu5CYCIQr9n6ZHV8Ko3m1UzH7Fx+/SZcfve
wJCaqo8LjyFngY9Bm2uW7ReDSYZ4GMaVB3sF4NShdWAx72E1kky84gY32AcwSC9zKb00dN2h3eIw
ekXCdsph4LFRqddIG/FfbQUCizzaRcQDr6+tFImRCvjjHYbEItSBFjYHH6oqyyFq+RF8VHeGS9TN
Rgnkn9PMGbXGi9iUAlPa9uyCkJY7BbWB6RmybCDDq2TfxvMNNFAfwSr2oCimTacZsTEXHqqP3WVg
uy84/2DKdYGLIxsCEDBEb500KfD/3Vlfs9R9Xq3D3JF4uHRy9Yj3ykRT9Yg4d014B3FiV92s1Eev
Gx34/IGtlmePe/s1esUdqDjuS+PvTEzg8SU/My5i8yndmQzmTbThG0bWUJ+QqPVMzM5AFBZfk33x
DL0kpmicriuQiTBRhXwsRC0mOB4KuGfrNJmxHo30t2JuinvYH6jYXwGm4a8k3n4X/n+iixpVBth6
dM251syQHcvSQpWCtNk4lBeM1OMBVab6fSkjq1EGNUDQSfo+DBSug06ldUnaOZkbpwUm1GqDT9sC
xXAyM2rku5C8dvya6oO5bQiYiBn0qmR6CasJO8xqq3xVtUNq1TEfUjs53EAKQ8525fy46UnXrWFp
3vi3UcbuQVjzUvb/O4uGGgAtjxfWicgVDAw6iNIFdsOvPdcxL6NuxS7UxI51ucBEPtXxxYIKm3uF
QkMdg+cJOKusOxLBgtnnMXHnEAWXuyTP/jj58rSKJJVO/ukHXvnKcVw87fVa4ApJqGwQQtIvrB97
OjbfbwMXit7D3mn+NdYibCmTNa9rWnZSi/Q4UcwH1XYpncrWpYPOlxKeufBnDMOD/ciirQTuM/0S
TwgnueSbUjlsaQLfZmXpjYko0x2hCeyYstafcfPAw2POyRMB2BsN3FKqX/yq0+TfQNa15N/L1WUV
CDrW9jsBuwX09raRG6LuSoxp73pLsqtK6Pv+x3l+rU04FEn3s2ZjD90yP387qXxiTLvcIHqmTh/K
6NnTte7Wd+aQplCrtSl9iuZlSyBUMxMhF5grSTbiYHOXH0osmFE+6MWQxuxjas2c/z84kKxrboJx
9vmYpRdVcSjFt968ptu+l6T+Wgv8/L07t+ic9gatx0KTyLs6VRTBPqmddLzwsOc+POGAboH5wDpI
foOyBunfG7ZdAF6fY9Ju6kOgP9R/JCW3btcJbOuyBlHk36xNRlVVasjtOgOiLmfw1tlAFD+6rRDv
LBIwY6JrIlC5YGrSwHMGNvSFsuCg/k8c8Zi7P1SggGNcc1MTx5A5FsnGu5p8Y4o0RyLHqLK2IDxu
QqbTh2+ADzvNQ6jCGHbUgx/lMpScdsyPJg3ZXaaPz3UCXO3JGZNLOYd4qLWzSOmxLJg49s5KIkDQ
AbdzgPirEx6H9n13T8Tpu931gAQ5YLTQCfjcamFAEzDpYiDh1nTEH69s37pTSoFyKhiOVzTQMp/j
1Kfb2bvmV63mRK7LJLbGHjCr5KICZfd+ljfNiQo99Q+PVd+YqkbuX3l+SrX6abbdA31M08rcNwJt
RLWHKVyMlZgbC/w891PSpWjC3CIuFAQ22YfbagK82SUlffqWXAPFuvL3hnLhUSma1LIBtfx1Q0kv
1Bnq15N+cs/yeM8isu94rRfNYsYf0ZfdTJlt6KL3iCCcW3KF9jweC7wEYwl/UdkgwWChwaFuf3pc
eFnudZ7bjLysOgzCPmVSRjLqrqkoI4a8j1yvfBF2QagsJm5w117swKq0sQWjSLZ1G9lYN6mdyidq
W23tf+PmpUz3fKg74+WqZ+yiA9yxVubzcAOu/t2S3uiflNT16p8lj329oQBkiXzv7pqWYox9uMgf
rOowgO+f60PFhfYcyT1DY03eaHNhQRpvUvUGX3/dbWoHQTdRMOClAkOl90fBu2WVjv/6c8Aj8iP4
Mx0bjPEEkQ2EI3XQIaUL/RC4qVeEkL2O3slrVOHxOJvJN5yPeNzWbUn9YOxFJtw4PQzcGWdW0FED
deku2nEOdXL3qGVS8kXHyd1aCRrkaiC7ZkcQcJ+cbk4IIeiQzbB7EwBSjQIzptvfihAHxdBiBU+Y
95WFArv+WdDjnqMgsXCceJZ1VdeVT0GhzUccCsr1eJvsPlYHupgEPjZMNpZ+lalX52OALexqG3C5
KLVXoRjxjTTq6GqkUBxTp/jMZgvzPzcNTjjaKtDXQm0FkVvF0X3F7Y5QM+P2MXM4Yf0ZXvQQPHgv
MtsoLs1kh1TvEF7D5cASrBavDjNhKceRxUysLq/7X0wQ0SL0nRD95aDdbcOSe5+24iX2d75LrvHj
gbRGXUgsdKJCfYJe1YvyxDv3FHo9sPACSBK5M6BJUisUBwVSFhjE+buXYbcQIifdygUPo1m8soDS
orJGYAKMCRzjZ494CxCSTdAGakPOLnr4yzCwwLV84zMS1vLrVb8HPqHt1KNHfqq65nHcn5/LMGjF
r7yba+Y/9z+dbrvSf17jwOq6NZGYL2tNLZkasA+eVNARfqp8sPDlIjPx6yn+Rq3npuGE/vjSlF8I
Y1ZyITJDmiisJhRmtXec015QXYEiBvS9OJYOKzp/6gs3sTtzYWO6AOK3etpWUV0m+RXapn/5j6J3
EfFPxEGWKKLShBijdo2/DlYAl/URP4gX3v0rD7FY3jh8exbEVhzZvlTcvEDe2Je4dX5gyVyHMmqT
sbMVRAz9qkWGjE1Xct5qof4Oj9wGf+twffUtXwqnWC8pDqwbF8GZ486920wCXY974c96BJIZmMO6
XjyHDgAD5Wp45jLJErkPYatkEM7Yi+iL+cnz3xFvBHZgJ9Npn5u29VuRPWGaInKoklMaFYAu+Ual
ck14fNHry0H+Qfn90FEGGPM0ciEa9Z/5JF+9szz70FsrEoGiaP/DNhyXWXs/JZW/fOmJwRiI8Ywf
jhfg7AyNu44b6MYUtHZYCUy+XpsMTnedg9YD4uxvrxVkB1FIuroRn+CMuvX9Txvs/8SeFxOIIkoD
BHSNFPMl7q6JDAv4co6Wgf7xU3QDUyr0jqW18hTHECzFgK4Ju9zxpDSSSuoRN/c2hSvJ/iJysjiO
cWd4xkc9Ikb19CcFXw5S+IvcWbfwNl9wXuvCnN8C4PKmfVJ0l9Ix2MqxdGvPGAFsR8hQsKScDfvv
BM/4tUqwPNE8R7RvNtk3gkDwXf3vRQ5R/0XXTQJFLJ+q5IfgGpO15nrttQAfEuX/h9PCeYqwYlAv
/l9SjITsydkWsiP8ulcFwVviLPq6zkAMNoUa21zuDNcvMr+F1wuGT9YsiecIL03c7G3dEk7GqrnZ
zKY4YAXPa/VPqkmoNGFAGKVe77ZYjPVclE22wGexWJBUp5tQyS5A70FuhzWWMlwyiYh+n5LHXzFC
WuSluDvNtUaDd4f01JR20+1rZ8cOS/Vq4r3Jw83OmYH/gyeVsiRe5o9uFAmAD8mMyZCsr+qoliYJ
FwMVKATYmOSFUZAgzLBfNa3d3w5i7ADn5cpJJXRVgqRqKEh9lpbKZeomihFqOpHb0O/jCKtfAIPJ
Voyf/SrgzJZTD8zx0INgJC8OIGjMgHjvevXdSYpjXbaiJB1rjhyUKwbT950bIrUprWe6eqLrRqhn
quuZ48BScRBzQ1dMBRvN039OpdNoSIkOk+UTBjvS+eNI6SEGWg9nTZ0QJKCV86C3UBzo9I9juiKQ
BjdhUdZQPOFYtT7JdHQk9ngbbgLRXSO4dARrBufG+7m+KVqAMjU+1nj8aDgJL2EoeMRDcx/rMaRS
wafX99SzBPE5pGmRbrfxx7Qa3LYxd5r1/DVEF2FDZb115R09XeEr8rFBn7GZ+lyopgu+deKIqU3q
yi1fxEnF8/FDqd/hWLbvz9VCA7cwUP2HHazoy2NLatqcA9+jq3nFOI/La74SmVQbyEt+pKCUNVkA
NDJ7lfUW4x1RahBu+0G2MpeWzEsS4dLI1R+d74hEKkhu5cTpw8hpb4kOeG2Y5ubRPy1+FK3noqOg
t2n2Gul5EjaVZruMJM0UHM8MvqGatc+NDSEovmUWJDypACyDs+adLPvCAoO5PwStqeJJFnJ5nYSM
qxYHrzwBeKFRXOklTGcl/hWagvftIDXeYufpRLHw9xTPEYc6VcAvPlhOO3hkr8V+rdEu60ir01Ud
wvWmMdi7JqDRIkWC3pg3XQzdrRvC6OYnf/D/7kxukM78TnckklO+kXyGHL9kU8cn9TaSluKQh8EE
1jYcW9r/Ohr/saoeApRx62FDKmufuB1Lxa6+gJjIWKCWhq7uPTenXLC6DUtdUSUUoiUCyhUvIFPq
YO9VA4xE1gP41f48WAGH1WZLs6wroDS3Pgppzkea6w4/tAtNobGh0XiHvrwnEvkntP9C+tDgQUT0
GecYh2AErbK/FlisqvU6GGHQDyCY7h4CoCuYh7JntpOBLYBw5zOuY3WGiUOgWeSBVNOgmbAK5I+j
tNveS6wow59fVcSniGgECocJNqmlzvZrpR+rxP8fLBSIpxrCTS7AIzTiIuvxTI3nuRvMF2dJQ8R4
AqAjjJ5TT2SUwQCprtgv1P+vqqxHvRSae4EtgYCAnXukG1JDc4DZUpZACT1XJhRvCFy7Dg0sCZoD
fryxsRaH1axfrf2Dt/nogbEnUlqQCvjNQXpKybgNn/CrU2G7E7I7EdCroaM040JLOOWxmX2InUig
8I5VFi0GJ18vUQCgxAvIvcZGz0CsykxrQ3RpXJzTRKUj//tIBIFF6fwcMoKvN4vggBIfz7/iy05b
oABzizWBuIY7X/cTtFKhmCUjEDWUyzCpWEeUuMRjaHDUTldWyQhVlJhz1Rd540Zn8Wp6ak+H0Sqi
T28ztThGQ2jvMK5IWKTt7XHieSVAjEQlJqa6pi/qaVslH7+8F4AvDzF4gv6Hf0qbEMkgop3TF7XJ
gkulxUXz69nzAdx4CgtjyXgV7gORmeoY+Pz4grGODYq08xdS+zAh08WbVJF1/hNTxiZhET0IQEvL
ilrIjLWvgBJsnGmmWqCbLBdFYGAx3VcWKNzT2qGVtKUvyyw+bElJ5MTD4txYHxEqoU6DIbNHSYn3
aTgM9GECTzkrCEMmUlZ5wD8GQTr8iznpUsFLZ3Y+dk6kLb1sIc9hzfkm+Hcv+5m1oeVocwotOZMz
PTFx/CyWkSwLZ9rmxZmdqQ422DpUH9OTl0KkZPap2klVJnM7cUqT1JchS8j8hRqDM+SEbGoLfQmG
RAmf+YfkAMoeEFC8FLKE9uV9EkxT63F8e6Kp5jfCm/JE82jyKv2ApJw3TDkVmdn08A/XWnEq4qTh
p9xtK3JgRu3rhQsdGxIDkLbrhLJCxdNZnljwmy4+zRjGBbgIEk4vsy0lMp57OjBaVuHsUqMujlfS
CqBJiqQ2DxIRIaIyWMIKgugaj6UI7IhCGylEpp1TudADRfOJGrXywuydDXOqXEwDNa63bYe4YU1B
t5lLfsXVwELZ1ZDs9e0AxLvzcaeQ07M3o7IYP6cd2qtv0ltd4MGuNz+rfgYZzXXD82YO8iL60ZPX
ZA3NWf5CKl7pqBE3B0zypTg4pcfzcM6TElB1927hRH3j6vyyVVXXpg9b44adyGzVqR28rws3zhyv
OGQZLag0CiIlETN7ewFZDI4Imqn3hRsRRB80L/7Fo/6JbgDQsoaqsg+yJ5r5W4CxzYl3hVYdJw9T
ttCGXBy16P6ozJeuygKLCVky7hSn34dfO4jw7Q2PTASCd469esh7fs+PMwLyjMoNgzps8zZHFmxO
ZV3ZNgXJ3p2gjuVkhTcWJsOwBrvofYjmH41q9D8zeFqqCfY3leipBQDY3xeuNfhq/LJVqbd18num
LvmIsdZEvr/iW5mh9V4YMCtDyvMn2gA2DpOKZcLLH7JQiZRVpmdrpJgWw2j9IdDnQ9XYVGyjOT4A
5sIStz4eL4ZikCqVqUReTOcrb60q/l4/Xlkl5YksM42neqMLySLuOQnc5KqMYxEJSa0IdoRZfP6Q
mztJ4a8rnl6MCkVBumEkrtQyAwKKJOjBvAxCIMVlPoXt8uM03PGZKjsQmBz5cjv5isULR9Yisrye
82+Hi9AuZ2E3RbDr3HynubsAqBhmZrjhOjUJSqCmZ9qgm9p4mBkg7zYyoUDXSX5Q4PWB8jarz8IM
lqt3nwZBVokmtHED/CGSlY5RqbbPa6c07MaGAa1630OGjFUqND+m5wcuLV0WJakCovxBhzt+sG2L
6akI1phSm4dN5G/vZzb6mFFInRrAQ4e0XP5tfKsZ7A/JG9LGWDZDsIWNOwiVo8owURs/rJ42IAPm
XbGKaY1hrZ8t7MdUDKauGYTopLeyI+ckv3YYXxHzik466HXbNe84ccmQiIeVYTOzbQGzPpQd5wna
4b0d4ceCQdoLxIcD+1s7YfHgUUEfhCONtH6rXpad2UKcmvVaUWRPKARXGsw1+230GnEsTpqmI3i5
UUqAirJb8QTlgYlElXmNQpEVPs5g5IFLxoFKl6JW8yCVLTOWv2BSN/NCsCsIxr95gJtDrLiMdVJu
u/4lq8aZu2SuwvCJW12CsWlVkpnLTxZZBNcQhmHYtW7+DW/Fy2V7OEH8zrugZE5PADwFyr4vPPwv
K/I+YUBAMPN03KDrT7jhKXv9qyfvvWVO292qTeigftRwI6vdmhHuldcqUl1TEErFMy+InVyJwPCV
NU1A9rHzLVdrI7PYztuGD3/Xy4hsGlzOGyGs3MQzO+KA3jajNJIdfe4q1NBkb5VA1yjKzRtlyKoI
cY8WUcwoQBVz/TK1dHu6b1UetpbZYLdyB7M8AiTwUBThOnw8BVkfYbuWLq2ZS8yO3rR8ehuZu5aD
dSdu0cAeS9SN/YVS8SJMG65X3wG4QEjJvO99jWQkG9OVnViXZIWPggq9oHwL2x8mvU7dLqneJxim
Juj6z5767wvhStsokE8+U45dNkASMK7HZKMu0klaljWHv+rDzWg6pMp3fkHxM/SIiB5ePWuoBihp
BRSjj0WT8Kj35N3tXjmnQZ8n3jtndHl8Ime5vCRjqgMar9u6vWQvf5efTr1tHWtSRJ6yMmBHqhHB
rLTEu7f1A5e5spY3odpDTvGxQEcklNqgTUs711RzclTXLRlsHj8TxeRSUSPA/NIQZ/Em4aMy/UbQ
Wf9EFzddsK3Cc6oUG3YVelGZB8z/zAJgUcRwg5miNSTpVnmuBtmEfIUT/08GryE2NGe2wAWZ239k
32oCrUMiOfCc2IrA3dXv1GYa+kl70UehRK91aTXvvQy6xjt77+Fy0V7QnfRczz+ihXZWAtXmUGAq
eKU/WGPp6DaxlE/vBj32KHO9DxZ6LU5WRMRa1mYUPW3vZ+ZA9uJQH0trTaSDPbpJLM4n6mvHk0AE
Npc3tNNOD5Q+dMca0tHBuzKeHpQxNCznDBKoDrrL4rp0PoXPuErhTbluogid6KveYw5mMBlK00nN
/XSo8ZtXMXT4Guv7PqBP/80OkgAuOBpGmq/7mW5oRbfSyob047A/Q3q3PkNZ9Lw6i/oSrBFHwjO6
43kij4P+PED33Q7bvW2FAsNkQBQSCPm6NFKJ4t67HCf5x4Ef3Tdyi2skNWk1zfrDsTl+9VwA/oBK
hXTaJs5wkzrOhPHbPN7s1fF6+d08D91SouRC2r/XbkzTirGULB6PSxS9DtbPZ585nGf9sxooPeur
CNKgOej+DHHvk41Kq5fOgS+adcJ5RHlT+P5UkLeZSULbYendFW8mgLvpzwgikvpgfYZiU4ZFIhMy
P0Qzgmksjo5yvdDO5FuK0ZfuBvOKSr0xpFvk4fkF/B3aGxKVL8tMwAbC0tS9QH/OPp/r6v5Icwwr
OGz4f7C6PDghk1diNeO7C/fTfRoeWPW0Tk9V93azbKGIdxa7+Q3vYGJ6SskJdmGu80r0oz4U+5sn
/luq7aI/PzLieFp9Y/yRGyoMGrrPorh/4WgDIXb43IrJugwjl1fuJvuZa0PuVGrInuxqqcntr3rh
1O0hjdUUv6eE8Smztu+IlDsyFAyH0c4ygeUB24OeUxUM+uI0bmYLWqGhQb5QRAyU6s4c6Xs24IMH
Onlha75pILKlrI9GnrzxBmzgQqS/idP70rHADPJ11wa6voW06G7X4jar2tbqN4mIgXhZLlBfH7Le
8fX0AqSW2lw7MCZaMnCeR432+sypp+JJvMGEJfOOm/ls6OVuWHyG/UMFNNTSbFiM+H4BQVX5oOaX
Uihhc5RHTlIrJL1rJFT3aUd5+nxHR+6aOnLea56jO3G9Y3gtlzGtb7tUpRiOH/5RiKCiPfPI1mH5
p/u4mXiUtHJbiZZGgF1lekCvqTfcGJ/yZVxkDVmwjh1BlaL+1J7EjYh+bMZi6ne0wbPbV8/KxMLf
Mdhv7DbKp30yGAhe+PRxLvgljzvJZT2j0Hl4edmck6iCTkMrxJJHq9ccihygwHzV24zQz3ur7w5g
DEGU2+b3Mp9iQwgeCI/R9F6/g5lYpMUTxB7pyt1Thi5vuQzVacj/hab9yfHqCrcKsiLWX3cGpQMQ
YPTiMFnYFwg+7ngTmm+cAqBrzU6gMsf0edHu4aKFwM7tEYb+XqAtLZ1lCm9XG+c05mTMn3wHs7al
2drLgrvYRUvG5Ly9JxGKtA/yDKh4RR4kJ2CliE9dxXDOXgnz1AX8FZJhK9Ec3nmLSBsRrWir3Bgn
ifmLLxcVixr9BuBbVd6W9pMShE7wyII4yQpiPQ48XUXa//xjPJjiVpw9roF2NzWYZg1P64ZUDo0E
hIBnbxsFCN+lq3SzQcDUfgVb+b3PkBc4dQOqOx4MSQY4QBMCcogt0bgxYwxUR/H2Jn/66oeOIsCV
q4kZRIAv+ddKBejI4l3yq68PhK8M7UvvAhfAon+d16hbV2MCjg/MOOQFZxQN9oCqaPW1Ym7DFrZR
GFDW6RFWZ0rqskKdszoTYTVI1F87mH+poo6WuHZinN+MtX7LRYzgguhBuEvKjIiB48fpZPCgDOVf
fNK4ZkrgtH09kO1QgGO1PTrTnzuYh4hn0N4QcwV7++6c/2XU/DzR2dVUtCoFsL7ZpTKLjah80tnw
E1JLNv+ON5Xeguq3mTtjlnAjnBEwncG3JBcz7TuQT+fMMZ5X+3newtRjYXA7+CSYWyT+A7Wl9ur4
u0GvhyIWX7rZp7lzddccjPUkfG/palrFspndD0yVGCCld+r36lxfYxmTL2u4YynP0AGgjzxt/RR5
1dnWPE6y+y7JcTaGXijiYhzOmmgsPd88XDsdaRIPx3bTLTqkRQ22hC02WG2AR4ztN/7A8jaAzIX+
p7+PGmzGCIQlaVT/DEOXRgX63wxkCFUEIkI5lYHXG8YkEWi1w3XEBHL+735f3pFY3WCli4TOBU+D
hEdQgFwyVxCnB32tlJAWy3oKtd4zRnyBlIWIsCuYx/VmmpFw0S/ObdvXRUdxGpHbIJpw+DG64ALw
+7ionc6CjEaGXxitsWMbFtZC6jpKeF5ZJLLQPduJTSF772zKzNHymPfBfVwEUY7DJs2DoKhDg+Se
+fQ01OAT8NpvRBtu3UTyC6uT/vJUzwI2lN/tkC1P5N7YXqHX/3i8vbo1pnTIkhAZ9hoN0bhl3+OQ
P5GTB4g0PSAvpArbLebuAyzYk9flgaDWU1a+ayJKzCMQ5p2Z6ERQa8/TSXnAS/Bqs1MR49rrbOCt
KJRVxXpuW8D0RGbdcpw/NkqjJQBEunTAYkhIsUDdeNNCaMazeQ5kg+P/ExU+UKOc4tvMKE59IFUS
RzFUVytXwVVxgkGJ/oVlR+BpaM7VzlwSEzq8jpddgTxVez/i4iMX+i4onPSBNSVbgc+5YxSgQJBj
i2jf6torDhv52bowZs+wa4n70xxn2AVaKw6HRWq3222mYlCFebUULNhtK0tfpoS/m76VkxIeLcO6
EIl1Xv6rfP42z6tpsdxY4Jo7QltFZsxu35biSKyAb0r9OktEFF4vQhOffnJepfe2GpeIVB8Sgc9E
5B8L17U5vnvV2dlmwzF/vzzZjW599QPFs4Nva34XFiTpOmXLib433ccMkptsFB361h4ufNT+Mp5a
zjNW6ZRwxytortVZAEpFEpja2m1z/Y+PrXEH3hrowl4WAejXmANGy0iR1FsqvDU5832+e7i4j0Yn
lSmwrF8NZZbODQcz11cvx6R0AZfsRLmRXzCmWJW2gvZji9nGVc/htDNnV5/fyFJ2hs12EspCSGOG
bMmR8N22q5VnZNHNSfHGjqdwZbLWnoaVluIZ7fdREaKOu92aE8zn6Lnw3xZtkfHo6q+ABbHwhYGt
sifs75oBpSO6JZ65MSNZZxmLxmwpHg525iJqW+HAebabNMw2yEVigfyf6TmVBAzLl4vXxwIruNvE
OrF5zTZKR47bZdH5+8Ge6mmWX7eMCBBF4ydXL1CufEyqRu8xNgjF37Xoc3l/kx/HVY48x3oBnIez
fPlEtJKO3tYgufq0t4RJLYJDxSzftlGgEcvoo7PWxqyJeUTmk4plEwXrYpB2wGSFv2EFik8v5K20
ULt6nhDCTIqkq7gL37aFDZjFd2s2cAcVNUwadVTnCKC/KOz+bjmg97dGX+oFCbq+lAb6wMTC5pOo
Aty7Nx0pC9eOoX2d621rG+thk8J2t19O+QwYOjoZ8AqQ2JfqM/D7aGBKP4EztFj0AS5IiiItbgU8
vX+jbpMkbDi/Xx2thmYaYIrfQ6akZCi0U0R2SVPrisP+/haOav1PMPBlICPKIIfE2JRrfurKVt0h
/nvZ1OGk1GbMdP35pVCLs4EaeU/QWI1VDgZzX/UyBKEL1Uvnka0Lbezrkm+dr3aTqiZbLdPLHHPz
RraVm5GBHgOOUE4asOmrNYAyM3cgbzgMLiw8cGsZGePdEu6MrKxP7GJBPcrg8y4GAJ5aI3ChIJT3
MrF4e9EpTYVJHmvtwC6AtupHvj5YiLa204+lFVKlVkY9UzSQfICFkd2TGNLBGLr22P8Y42Q/yISE
3cMWpXB7xcKzcBp/16Ep5FyR2+cxi1jZ7xe099gyiAyOZxzeGCMaSJk0oq4/2/iVLwvjGYnSSrjm
kGAyc7t8UIAh8HpO3Ez60ygZay2gZI9amwI9aiSGIKwkVMwuidXOsDjxMV9zkRPVw0gXeyXVBRnV
24b9XOxglgxm8GDlLKypXAFCE66Ljf8AHHjubtBKBt2zwOFqKH7vur9VFD0JdQKd9Z654UsMtAF0
ar7y6DbQGvkI527t/UzbNMrCZzDfGAOoAGBQ4rNd1hXWnYfjQt0Mdke9f7A5gtwPo9cOD0D9uzX/
WnIdyqSKkTSJDEzxrqGbXHvyKzc84mdbdVIyBVdbKsgurVcJ81JrY7K86Ub4UqdqrSL7vqSLt/Mc
x614/AX+7IbiNVnETOnC+5LJgHatpQorDIJkEcUn29npdgDdtW45MLn6rE0TUil+WyJk0cCWj4z5
60NsqTKt2Fvxes1uesPJIvmqzx1GmiWY3LHLx15MWB5XNZlrk4vSWYqbRuKvFwWTlIp/HNa5gdg8
j7jZCqUa71pRoNZn7xrziNN5V8LwmjwXds6iCAC+dodoSMCipXH2ARyjFpq9XJffdRptYI3UJdCK
Hy7q5kL4/DBs7LhGezq7j7y4OjBheyQI16dzdcnpXJp05FGvvBWSbCk1Wgl4nf0otR+N5ey7YZbg
hKDExXszBJnHNIpddNt3mRdhITYQhmvaLXaUDeIRES7Zqk8bvP46k1B0E7DD+G3QU4KA5dd6tUP6
vT+UAtQiKY8EnPAqCgNOtXTU3+/GFs+CiDj6viORMEo61auT0wQNgLpvHCjBJofvOBnwCqJs4CBF
LtG95f+4vDRf2JgkayGelGg74+TO4Wzv8f/LhO7/bQKWTVUOFhuZaxKgBXrM5tu6eTpfGrDCjgDG
Jqj41Kku//XpFvCFyngfFoQrP7K8eWnS1XBDM8xLLFAcjgMP4joCzwNIgdDMzw8ARVkEB1MIOYyY
L/lQnPAZmBjraXkNJwGpin17dhsAg/ZhC4ZDJU5pY24jKFLGJfAXoUYOnpH0czfqS3sGjAAUdLo0
ZFtHnMnOpwmpFdCf8s6oDjtF1tViyUWZwNvwFx7yzc6ltBA3wSCXghO1PRCjgAmo8ZXczHxWXs1H
Z93GjvpYNWezKYq7MwgGjwxYTesCnUmz+bYLbkqoMPn8h2nNiYEdiOpRJFGaFtREx9RPEQSOyMYD
hot5ocn6j4UZjqjHv24Gel2GDgO9gT63aheJ7mE5iHWa7n7jusduAdniokfOpWrWevvQbk0hBe6l
LLeeSdUcSudvOYs8pdXApEf7KpKVAtqJm2eBAI5l0rGmd0XEE+tNg1IRDtAJ2j+NvKveVgM5cjHG
1aYaUHjOH7jiFCgl6gV68k6Y6ylsdbxjMH1ztgB16Ec4ZavJW3frmqMhuXbuF9dxy6hEiDU0euXN
EHVUCxCcuoEoGr7YjKNRqMoPFhtYMJ9dCa9m2duQ1QP8/F56szQ4UpSqsH6b4PbKYgu03JEqgbMQ
q/L3QZIY4LROBNHL9QOKs5wsll/YMkXSJmzCMHin8alneaE91TbEYzRmIBOGsZZv5foCa4nMM3Mj
lBJFx/uWSXPvaLalG5G5dkERgefUQs9q73wGrhOPxJPVDfBDYkmPFdiVuA7KV64diB+qBY7Q4+6K
eB9o3NqpZ/hfZoTapWtJOwtcE6hNe0Cr9EHAxACI4uOtB5NcOx/iTCtMn0VPBAXFa7HFLIpEvmSi
9NdG1u4vi+klYKXRJyuBLmzhkxaxwXfVymh2akc0ddfj72D13w1VKyU4JhwpxH+ckmI9FvwUsrPA
8RxjT4cpOiUiTWUG+fkjVfUk+AL2Qpf2EMwIY8ZQiaSnygaG7p1oKoPVunr1FeV4azp+GEXxkLHn
6vwGswrsVYKWnmFeVg4lDOUTEvvNXPPVDVBRRIUY7TpihbiRziz9e7ObnucKCeptFJWLZUjqNRV3
mnh+9vnkOTL0teb5zR7btQvLrjkzGHZPjmUky3vI63ylJKbs2eZnwKGG/hcRl7QtWjolskDTRPaD
y1ScT1ns3ZfdmzCE3XVobmBMkPAkg59VKfVh69i7/0zg48JrgqPtqrPMq0nAG7NAzE4f1szjnZaA
CG2WAgm9NBIzjf1a2cj6l7lWliQwGScUER03kBu7JX1+rRVyq2xh5bOC6h2MkFfrapkWZbQo5kVz
7IxMTjRLrTVOMn/5pN8FcBs39fb7ZL/83LmbNoBxQlm5BXyUjWnyv85iOFx76zsBN7RE//SfNL++
SeExmBVOpVp6LMCjr+gc/0jTJMC/WXUAB+ARQQmT4Zi6SjPA9ORsP9GNSC+mQSFI8d8Wo1G1eHFV
5ipJYeIj0PYcK/VuJfeVhQykz52bAMyFJem4/UsP91EOItV3gMcxf6x4oP4maEUikoJ8Z+xKy8RO
Fl2bcnzgbyonjXcLMJIe51vQjqHze4gLpe1OJwm4TeLxD9JgLIgQ+edXKecn9eVnK9KrkAWvEb5E
k4ePczKsKSRjpvg8jITA63B+33/TjIKWb1ytj+mIenejnC/zEUR3HTAivD1Ck9qRC6Y5ZXKYjHxN
oEHOvxvqGthAopW8K1xmkfyh56dNu9PWSLtfqrizKkQXLgUuCrtkocVxbM9cDYknTGYRlBN8ak33
gW9X2HNqQzqjz5fyanDgaSSMoFgwvgBmRzuYkcWZjYliR4F+hJsGai4q7rqOs/Ux8ZWchruzMUZd
ndsfITSl5ILDI3HFqUKFhF1dCLRn6O6nLj3wHQHjiGi2gMQHvqgbvzGVyB51zQj8Eluo09j5jd/d
egIPn91OLuKtEOiuFTNJx78tX1LXNRMwUTFtwCYtOueFvghtweA9jAbm8JVpt3XOPPM7msvb5Dof
wuGhEmNwGFqaZKy8Jh9uQVSNx+fllVLRDdjecqIULqXYgO5bFlfjT81LbdZgtPM49B4HBqTse7f8
5xuJPeKRCOyOc6+k4FKRf/n7Raqy4EDr/lTGJxMtzuXiUA2Mc7lGv0TggrwgKTfeMgLy3cqkBLTv
l1X6eovN2DvSOIVYYu4eENEBfn1NJIuvKtvoiOHYyTZ9ipbQTVYr9Sl01RWN7mqh6RrMzHEvg7s5
ehWMwWaVdjdCmYY5FhJHb/eEueZomvgPqPkt49t0AsiYYMsrnW5lUP/aYPs4tO9gI1eTU9suI0UI
G04zzM6z8u/RpSg4X+JIpAgmXnDkgW1gWq0rKDZonWbNwp9/zmJw/eAOw+r1TMjxe1idGW8W/m9p
KRfOooOgia0BW/JoN7YP5izSw/yWhLbPoFeSkEMCj570SsA8ZDH2XKxanFaDWU5y7x6Ks/RtnugK
Khsahk7h/gK8QtDwO65YN5vFCIt7xlGAGzq8Z/EYxIvM3A7FXRzwB4hbO4mRqT6coqEp1x2tcBr2
SzIlpHQtxAlGvOAEHX78vSOT76JfIm4gV8Ea/Hn2Twu8dD8b6CbB8N63efUxBksW8/Rdl8nhPs81
UnOfHwQRHgbpc5rDvG7UWDJo3OwsOUSbxJyVw+hFINs7deiRlF0NMpXef3r6YOOZ93emE3RQM+nY
jDu8/8HEyjnDvXnn+5BDvxK/dUdm54XspnVfbO6gbHQhzEBylpj8fq0oAbm4z+KeJ1bfz3xCofkM
XAeoJViSCmQTi4koAJE3ZHJCgHXqFrXQSkfLvkodGHDbEDhyP7ZAd6BBdS8ezL785RDf6rNc/OCe
j0yOjQq3SWtp7Btj3Kg2DvWNbLSjUWyp1UI5ZD9oGygg8e8ekFQ8ZFCQyr50TWBmfUZdN0PQaJN1
OC36VgUokbIDs6tZ++8p1aQLdYo0I+MyolKG1cQhvroKpqOjtXURpV/kUtDSJeDn3Mz1Rg6Dqghg
jqOoc0MLi8OXRMUMUCUk/k0fhYjcxv7XicUvEH/Vzc3JDG1hxeyJxs8FSwJIxMtRvKtB1U4EbeSz
4L1kW9zwH+VksCfafhw8Upsg+/uMkQX7pQ9d6Wg2Pv+BoapJ3gbiEz+ToFMhV9y5XCMsvZ83Vv23
P3X1krIG7KKxxr5kJ1DqzTNi+UZUQuEtGpVAltabMYKUxuvPdoVCvTPUIGP4y80s/RUKL/HpwgJQ
3pWzR7RXTJYGMZWqGO5jlCviRLIzylBcCDeaeHUJYdq8eV3GfFkcqkZ6UBX0S06E6ESkseYjfrdB
xmkuX6mbTLuBtr8JYantvyiQ0MNAwcjk5JSTM3M3GBwqEk01hB9xnZkAH95XJPAHd7jIxiHzkDJL
0upqoBtNwUoIopZE1uQLlnYBoJc/BcRwmJl+qBzabvMpJz9Tlyp2gor2xmo4vUZUC3p2nHAcdaHz
ZGqkckr3XzFBpjcYfutARM/BdK9ZJelerl3AmD5494+Mmqgy5sTiPGItqXRJ7zj3Gy4s9GmsdKMV
hfunu6k5+OmxqhzjxYNTsJGmoSLPjix+KNgPJ1jGaGUX95TqApT7tS5myyZbvOKF3YVwhIOVzwck
TOqAafOpaRArX+fwz85zj/EXeMEIFvmaXQKvot34fH34WJsAS61pk3WUfA/TvabT/ThN3khXHO5N
QjGonDgPW0M6jMOGOGXH5aYidenjfj69pTHhaXjjWoaa238xvXbWoxoYxjbPbFRa6rjznZs2iw0B
HjBE4wPKoxrxr9Ujhc5QG27BFxXdI8oIZInozjMsrGpU2zvTZmWJD2GQQduInWcv7NCrInCa/q9U
AWfeL4olbOWi9Bu0wQzwf3ePIk5rh6+29bAdCdO9zzUilNIlwTK4SstrpIfOzlcxUvTyVgkBOACb
+i9y1JWiSiieWeeSpb1KTpBnH3VmL0J6fdSQD0HUsUU5PXJ3IFGl01qxE3A14UVRCdK6kBoHornO
WnW94W/HefAmWQOpggNaUiUv4Zt/UPcLN5UeWOUtg5rRbhHvhBgdFIHQEQrzbfUnklLApB1Jg2tJ
J5NB42dqnlr3n5mJ46Wo6fyPCDlTUqzU47tZ1cm4cjBtjeVyU8dt2nfEDVvSrvyL2BP0TGRPcRo1
XX1jtJCQQEJe9QzEiFLBznJ17iFILQjiuVksCwPxd+vLUVWITjqqiRHxIL+tT1wKZlHoj/xFr7Fe
XweYCc9djFfwAAVf9CgYFlvmexGWryWjt2dbqqElKHBHXM963cDbW1gMJUrjOMJVadgKVsPRdzyU
wXlVV4i0RyL2pU5WIJtNU7xO8lHKFEBhwnDSQsgyiXluLfVhHdDDD4ERLePXO1WkWPcdYn2ZecRR
GkgdB2eBGh+q1DKVgy7UuG2wbHkESmLIVCr48fTY0TGx3E4wyOkXIwmMF6fkhhCRaEMtNzqLQVXb
tt1kKNbQi265Pv1guHQaisD5A2FWVGzy2ctQmgltQFuUiTHv5ABAA5DCw/shH8t7WE0MmaRPGxP8
fg51gsVhI970kIA/CS5yQQDx+ilzNUQBkMNMCCs/1MQWkGfjqQeVMtbvkzhQofecGQc6bL8fG7D0
rOYr1CSEcHnC23MvHLwbTfd9tnlriCUfWYKjvBLnoHGPrC83gFVtfTCKla6x/r+ZvbiMc2QgIRaq
xATj6mZDa4RtBpkyNNYI4aAbQfjtGyK0cmIpC7NJvpjW+ouH6SPIO/s9SEf+Asc8Poo/GzRi6beN
cqJ5cd0nfyBY5WsY3rW7263U7wEANjNk+IsUYtJJfTb9+qpbDYov5KPkj0YUGncLgrVkX7qsghY7
SKaJBEAq7yYABwS7lcAMerR8SJp76vWEsLhFHcjet7I+DQivJGbbhrwFt+9NV6bcLinl9M2fL3Vv
Z7cw5b3W0abnleQcuXLgnTEkjR19aZGjQyrpcaQY/eyVfoS2zzNc8PZvu5o+mb3zHc76AWBBtlrA
9Iz+5BlqmpmyXHbUiM2hAWXTF/4946unr0m7qL0b0YnhfaJltoEsyXFUMOfdN8oH8R/cwjr60SoU
B5ju6h4PgmD+fO9n96NC0T95QgCrIuli3dD7mwmXJd7MAy6sY3awOHk5YqgoUBqavfcIfYSTA6ty
5qG2RLjiQiDHSj2z+hwjg1XbObwE0T36KrHdSc6FXUE6OWe7KJyUsX0ZpxCv+YESOQO8iiquD6JW
ijOtffIRgbHszJWSSnFN1z4Utky/vpOFJb8/Kqy9ObuE2ynYt1X8Mj5D4v+Q6A79wj7F2+PMm+Jq
bAnCO1sqC7qF/ZB8uLk4u/6q17jy3dbtAka1haZaL8JLZ19s2Uo6oRwF6P5vI4lAW4Vjhht/w6bw
oT/fuHW0DU88ncob02qhYnfTjAoTtt1Tx8Qk5R7A64PzEVGnVkPIXvDJ6i6pXpQohNdrJrAu+npD
4bOwoNe3vxI7jhL11zG4Oq804jdNwM4a3pm1JVgPxGguBJAIaUICuJKiKXBn4KItyBkOVkB89sr0
518g3ADgnxfCRHvXTzyIRzp7MBhLgUb3NkSFgkSHuYhJ5ijBSIqoQfurIR3AxOi3lH5l3RB+RDxE
f4fljyWTRZuoZ4i5UurVn7Uk6rra6m7BIKF0ncqJOAeA0nhIWAxISsboa8zVy50s0zb+DkadXATM
J1ZQIoW49Z+10TRl7vefcn25YYCgqoYJp/BZiS5plZMM1r8IUReKja/i+w5upZN0wK75+BhO3jZw
SlNqfDSix/7MrG68aCqYVrcxi1wSZk9LyMLeMpJR4fLf/VtDf6jSXn9QHpkeXXX+MHL1L9yaqLgN
8fq4+qKVFmsIc7nNQD1YgGWFnWnBvYnPVt/cnLQykBLfmZgdbyj1eXY443bn4uOv01Pf4Pls5CBA
O8gElZPgDf88c+l1Njp5Y0Y2P1eyoRHZoPp4pbRLI314OKpEO8IpZVi/OoHFJr+RMlH3NzQF3lcK
eXxw1W0w68L1r4vG7k4GqTQH+bS6NNcsofCIjijJzRGsrpOevmlMabA09h+ouxWR4RV4bSq7oPkX
2h3YI8HmvJhMsSnztBbiCczgRxhpqRFaMG1wtBpaMFJyO+IJjFnfksUK2M0eapESEc6kLa9LIV+1
bfjyGVZoFCPQxB9aExdvAx0cbI2zLvd3NPdKiZ9P8ix7oYOU8VzCNgx3tIXFwE3q57OiDC2ohFuH
EknzoVqqdgeGTeY2tbs4CCAqxJqca+Ly3BDLafvwIuIHq9V04xmRtVT+uNgpy2DaUOz6aT60ll5N
WxQmayURI3h98V1rNJB8PyZHjNTlglUOjdKDBi9S9mMgxC0frrpy+SeqRYfqVMevlGCljDOGwFFO
P87qrqkVzNXoJgX1IVAh61EDKTIFsqtaWV3tZuq2bilxs9tabwr/IZRVUYVhxsebAaR6s1iOWSAc
l4AuYhCJJjBVaDvWJn5U6xkcSpFvdEDsz7MBvBhyulW1UNoTTXoEvo26y613zPvYMI60UsLYSPgR
Jk0JG1nurRQIxp7gZqmbT2fVmCqfITBSd76rz5R7w/5lk2hPCZv3bUBn629PUcZm2dMCbf5kxrZf
sVUPFG3g7g+qzmXpTOappoq9SWYJD+GdSnKKOIrjK1831tsekKhe8JFIrtOF/fQsVX2tPXuHtvlm
bLjnn9QkGr0fdDYuyQ5phw3rTIe59lQii+JqCxFRgTu6dfchHbiNe/12CVDqvaMrXdkkwQ+VG3Av
kOmqifQeYVi1rQG1NlfTsFWF+vlLK3ftIJQKSbRxfljVaYdK24F7ulq+zrc8pL+ZD9n3A0QKdY4V
XKv0sUZTEp8HtngZsx+XFWBKRNfGC+UuXbvo4hfi0H30vsldVV2mrwXlddgiOFZd/Y1wUPsS/LgX
jpyrAIYjnFuOCcTDHTnREfmOd596vsd3Yvd+HJ6jXikhD7R+yMFdTFeO5HE9FKS0tAj/1i9t93FD
yHayJyVXjyd9PDmCTVpWHUuHpnyvAkyUv9891TGM7aABTgi66xl3g+0W+ox9R65xfDj8m1gMr5Hw
KC9q3O4nP8RvBEahZDAsn5Ww1RvgVt9O071uihpPSY67zYPC5Vjfxo8gWkmpOS+Sz4dKJI5S4tmI
lSU4G3bLL16Pq5qjsJYGqXNX36WAxiG8FjKA0H5tEQw6PqEdkLrLu6iZ+luTfuUrkeqJdF4XmI+0
AkoqqsDklkw3monA185kj6BeragUNrgxi/lW5DKAGP/iNn0iG4HVlfpzNtwRAdeB7Z2mvYP7CCKY
hp7+YrGrLnXI/sYvh3FHc+su5g05Pl35B/E6pIHKrvol7GQoVfT7Lr4zd/G4Y7w+TeIXgCCSyCAe
1+UtcYXv70ohM0gBl0HRuGzCmCadwHqjCOQKXu3tSAMQKnLgfIrJKSUupXJW4DkdVDOmKciqYEuV
NxSwOEP6dY0K5rb0kypWL+ZdIUBrumU3GJcCqb2EkL6b1lydE0ql4WPSoDZ2tkqoSvYj69ECVl9h
sOMvkqJvD4hUx+gODwWsjAdrvDtcEmlXfpY9G0+uDu07SYIn4hRJR0xJNHl+i0FU1X+nw8zOml2j
IdrP2c04hjndcKS7IZVm/UFotNFTUhcGIYd+VQEHYteAw5BOFtiOQFAqjAxYC2X4JgsVfd9dGhkX
hzr7bbCxumXL3vY1uumuB5zApJxL2Ct1KliQuHMJggJxZw7IZBz342tsBG9VHZnyoWufVU75JAZJ
0re/5JQzoqpGpdURpoG+tFrV6vzvG9nOUFOQROYtwPgqzaluMDAUqbfalVaF3o0aWB1zVR2gFKuz
jvrbm8FFLJJD0F5qw+cX1o2Gga8UOfulIkBKC4s9xrlQnRBiEQAJyBfVua8Yjw+E6KhAWXsdoj1W
sN+1qD+1WgFxDBh/cTCY0dOe4yQ1qklRXhI9zLQvxA7TvVf8oKaePgPJxA2O0NGitglUMlhk8krQ
FJPzc1G1SAOTcIBZHLCdRKb6VLhhoRIRNvgeMid2d2/TUwzpHqrvmsV9bawGNwAgGBdIaSmf2Q1A
0XrFwsND7o1A4FDUGCkPzjafbKXbtvfksNaJdJxMa9GKII0jMqfGFLJuKGwXJb1hyGgJ5Dy83sVu
tpx2QcqRarnJTtbskEKXN67DihwILuQMd6Q2uzdM99UX4ZUeA0oqM+DErGlox1LhnLQvbBYtbV4s
OqVyTkQSJrQhHFrWdxndI8u24fr6Agp85xiDR4CSRpe1Ku0h3lrFlro8qSmbZjRK73Kf/ygjsjmL
zrOJ2wo7gaxuo2Lt9ot2utl2E3SuCwVUIXL5FLmj5sox2Zv82/7yJ5Yk4ZQRNDq/LgNPqV7ubU1U
q26UyG8Hc0VI/qEpQF8eAYj36mUtTMm4DMKLFH7B1gIHWOS0B4uACbJCrDTyzh+4VFm4Q/feJfFv
0DrUlKJnIuC8lyKrGBTm4WmoormmQ653cH9/MVpq4kaZ2Qt7aisffmpijcQ1K/qyxqNgTtgMValo
/FEMlrOpPxKxHYPJ8Dm+VfGl4tJMwJYqpjPNy3DRSQ9PNUsEecu7WfbUH7q6kKLTnFwUv5SzpA51
Bn8OgE/ypMwn9aC1We3XUrIdyRTxk531B2mhdUnDKAx197yVgtmftZ8gxEn3ogopCyLxFxecfYXm
UfwxKV/rNSbODD6NSahCqJ0o+kNW6dtK0l9lnQfvlfL6UndAWB3GV1kF4ILfVN9MAuV4ipogwlBM
CgjxnGKDC30FkXZNmS4Y978zu4um2P4+FM5EsGqgBglANqMZg6mq03vIHcDg2WG/VxTWH+FNZW7T
/PBi9JAkx/a9VpjHr/Jk1pBCuLsTkfHiSH37iyvAxTI/I0nj0aZoK6LV840Nwr9uKLurqjfRQvi9
Htv42Sg+sc/zlnJGmlk5FKC6SgG8f3YvfsywiZs4Qi73fGa8DfFrUxufSdLUdVzgrBikyBjDnlZx
5e+9H66DauKLbDQIctS/WpydbNq/aMatkTiC0lEQMzLB2hIg3mQ6iychqFHKNO6O9i5oPrs9kRfN
NjesWGYUHD9/XQEy13vqCZ45425tVL6V5RN6TDL/T3blXDNZ53jOjsFPk/VNctYwSojPTTAmOe2p
Cly1X0oAdLxnF7CDq6ZUQ5OGn+Agid+wO6MoL6nF05kD2YPLASpOm1yiQUamj/F/W6I/myzwEivc
N6g3M0wyjFqHBVarxAY7AUZHQrMAa3TVjjD69U8JTr63N3nbEXpV+q7ixVbF55UWUz0GOdToT2FE
Wyd63CCizxawGDhTsvRTZw9/vfMyk2qCM9xG+nklnM4a91h99xEiVF6FeBn0GqMOVUKMLLBbzjGi
C9oR/jqXvfXRL7LJo+JnzDl24/UDDlGSKDzGqU4x4kRNLolj3FVrV6agamVpybKd9+X3xGygHCTr
kTvhVUMR3dSM47H2V9lzckLul0U8LNmEblwP6T+88JULcSD836UGQOGmCkoUYiOV18y6VaONSPtj
XVkxqatjhoJRQtY1T+HFRuFrl3X9pJzuAciWj5isyeFFasIyP9HR9oc/1CQ8h6EZmuuBic2g+5ZS
TjpuMnZkma3P1J3spo3vjGHQ6dMF8sLrqTZlRQeQn1gEj9o/NV6u5XNBqAyBXeLq/6WGOJ3hxp/G
5cQ15W2HzPSRkJdpzFvrNs2QMGvOhCFa17A/97MnSojjW7h7Bq5DufHIpjpp5iImCB0kSziVUWJq
V3cHhAHouk3z0K0iXUcSlB6Bs/MZiub/3xqy2mE2isBp1R5FZoAcFcXb1G9lYQrmnUM22M6GzzeB
tSNZug2lqlw8zdsYG36KJs14S8gUucx4kmoJq/0ONmZpA5DFO9y2Qv+CnolbQCIPmjAhwnWK7Avl
P1Am4/B/b3dOVp22rFGgV1INsNokYY9vUuYvgAX1H76QnnyceG9zJU81rXEPs4QxiDWu+gZgHfJA
6+OWXsR3h1nhmLUOuAZwYFGSbPOA6q3pPlPBVz0QH+l7F3V5zTu9Z6yDfwNghm41IY7LWuL7zKlq
E7SJ1e6ScOlh2FESyKNk4S5DrSwC97NogyWvdy497cKgRv7vYboJtQhcjJ7mbLJ+en2KNbODsqhC
y3Yu3oG+viuxDIYnMb62hmbF5NxF5izIy2BOEj1XqASoZHHMFzmbm5Iv+nvfbFl8MMNp66u7ZJY5
N3pUIF9mbmyBargrvks07YOBAzEcEpNlAkrY/I5hVUtSPEXUG8uVVtHCtDe4cSIsFP4NPjYPLK2P
eC+GB5Km/EnidWiLQCfqm9TFD+QQGXf0NaG/58Vc2xg5bpG6RuaiNwarEG3o6hgrZHXrH3tTuGhr
V0+nBburREJ/b+rbl1RUKXiZwF6vEtFaKiBhhLCSWqmHvvt+GdgmZBUBmuPtVtJfg0Q3iYPFj1gG
E8C9HYtwLQ2ZblS+tyQneieBgr8J8Z5FUSclP1PIrrPC6RpSOQ6Mg3VpMdt2M4R7a9kdNaYdAa7F
0WLjw/pdLnjFBJ5E5vVdsE7LIe9Ypix1+HogUm9BRVqnGZaD8uKUZRYIbRzvnyb0nQEV8rG+0Dt+
7ZXVxi4G0frx8ZndrN0oFGh299eii5E5nc9aw+Je26i6Ezah1yKuIwwaTIArJQaHizyRES/LPL9w
W19PkzZPVdO5Wl/wc2jZljgI3iLdyJclcAm0YLCPKZj5vaUPYGdZYcOcHToatxYvu3UUflH69M0w
I9nI7HFzI/PDiAd4hjKcBi28JEJ+zBtnKRm75Qkwp0hUdTEA5krPwvlbOIqumY3U01nFGLAWNv/A
FUCeOIIpNjZSJSfBJEcE7cA8ZnylEwkME4DXKUZwtyPmUBFLJ+KUqLIDsTaJYZL+ARMZ7tiMwRqM
9gPo22ZrzXJh5JIcQxN0LE2f6A8fzPJ+kTY8A9PDeeB5leDZZx06+xj71lbwl2xGyLESQSsj8xt3
SOTdVTk3IJsB4R4Z7bXBLt4d87ub7U04QFMIu9G0q7WTH9+a5o9PxEDF1/Cehe2zhQ1efsyw8/IT
A9H8LjjPPa2DT46asm8RonUI0q3lEqge9y9t7pZjouuouYiviGyxIPEDe5j7Lmu5VGiAa/W7DlsZ
vnY1sIDe6n9cx0ua420LgSELR28YvcIRXBJwx2JC4235Ee4vZedC0RYiVaCfEFfcOqCSLZPzYO6B
xhnfOnZ4q+UAt0XY6LhdKH+tSActrd5Feid+JlGpHGnGaNKCADmXZe+PLBedpckS3uBbJvF84KGP
s1LKKg3K8Ubt096dXYzMyTm4igS5KCu2Es1vPj9xksmQf52qI7FzRHetJbhkvU4+z5yKVVJd9MHi
5HPEoexheWzeHDV8UN4itS+BOgcXDEXwl+3TADMdtIfwO0ahZkdOsoBi+WXUgLK8ltEXI9NFPsNU
u32yjJGs2IJz8ETUYpJdrk1zyFUsS9q4gRwZV2qRVtHUBkra1FDvrSRxZV/T9us4l0wIHmPuSf3J
4mGN+28eUFrzBdhazw6QiJ2qgUkoOlWe4tyGSHL8jS+OX8oHIeAfVKdSXmwPRlgOFxdV2eBWj3wK
efNl9LTTVwWBPeuCF41ZCCzoM+ytqtz72X4cjJjcxX/J36KkCXvoCrbq2NIN79SNDlgI2YRKEIDW
Xxhg36eZDD6TKNkGeuB+Rz+C8UI3gPEMaUpPa527Zsy1Ygln6FovVZ+myesX9OqxsAhEqWi8xt5s
w+RDgByrH5ORPB2DJ9ZhVbb+L8w0ph37Vk8B6WkZX66XyBaO3wiPy9yEBpYepO0BNmSnM2nUJB/D
Bu9oTFFPRPLXCjplNkXteS3zZ0FGs5u8rgHOaZ4VFSBsm02svfSDP29p+SJ0lxEDaXJVr167+pmp
ZiTc7gS/ptdGsr5SbnQJmx8uXYPhKLbyhNpQuZGY551/GSdQG7pV6pkxCx6bSNHG2y7a4UqCEHKA
OvpS98U3QTOFwzzknER6SJBaApqbwRe77IBT0PZmHzmSZ1T0Qmu4RtTHoLhC1JwrZH2Nona/ApEb
hUHntg5xICihvh8DREPDseLgSt4TzeduhlpAtLrdkFRs24LIXc8sueFuSHek7FQkeVwuP5H/Q3bv
9dyCxostCMkJpEZFGwGvzicU1z4UwRecF5AtqJMmSjdgvAk3U0F/LY1BNkEWQNMj/lL8gB2pCcwx
2IA9Yd1TPNTEnmtfCspAM55OZB9DZHFkVw9mJoLU/5XxX9bCUSjuHTa+gjuyrgiz2IEMo6vGcENr
SLSGZHR1XqcbwO9fvLjRTUiDTr0Y4CZG0+7ZcMl8dLA7aT841itC7R7+Lj0x+4mbcDzOIn93mVbA
vIINLQwb54C8clGrLGJIaLC/xwEEkRBK0VxZdqbSvAILfMfSlS352x3622rLAZX9GmjhLNx2qzOX
igAwtMKO8OMG920OU3Pw3Yb0s+oH7/x94fkx3Ng3v7OhIgfevRr95Jzw8rGE0PGW23948/CsrK00
5JHjR5o+FeXPb5FrTgWSv7lPK3OzJlma1dtE6kdjBzY2ALFcwjPsCw57XAYdQrHZiz83Qd7kpZ6B
ywdM4Kly8rjcXQ+OCXHUmYWCna4h/AuM1DCBSKH37p7Wja2uRlNSg0QMVuFU10h3SyhqHghkQS0n
Q2SZ82goAqupEFaBzr6xzuUv2kfkTVK5l283ItP6UmJbwYiG6Mxv5WupGl2vE+ll1AePdn/Aw/Ai
mpp32t6B20hpOuDnWo3UGag+8k7vebBi+5nAog+c0U1v3kViWrEzB7NuRF0ua7au6i8QCJemJ+fy
ahp0/xY/Ikkl3vsowAbzYklnnX9q/ji2NS8gPXDNdbhy4yfsfVANRnL7xeDDjqq9DiOylVXl9xO2
TntPGHjpp6vbbBVZjIq0/K2d66qAdsNTt0Y+0q0qX+Jz3UXApfC+0UDDbG/vvUBvI8X0BNbQ1tA+
CqHT98OMdzjUl4C1Tlr/9FTXLBeMdKL50tGJopYCSmRcW2fmkYa0KrBA/KZWWQp3BacTuNVobG/G
wD/9oGkdyr7apKRiKxL8DcVppj09+WoAKSJBybwlzvSHKPkORbvC/vaslhCkH63MQKNA+5eNR3Md
Vi61Tyij5Q6k/tjRQ7M4Ap7WJuCMc358uN1JAhFSUZAfEHwzDjhL80VbUAdqNabDTMhQlK7qTey3
ejwcPaFbbL/u1vNk4DL9iZxp74sWUd6ymRShNYDT8BW8hHORuI4hzSeCB/VbXSjfCJJ8CZBESTLM
7iRoy9vRz4Eu2zrsggISD5L7DVmbFhiB5yZsyEMYLtXLBdxRxKa9V1eSqoa6VFriXcc10pYiEsG0
e1D3IQjlcPVQjXx4vGHW7qiDomM7AMr1ZS2e90oNrCUUl6lyVSZPTab49+bpS4vlWg6y+xbOydzA
Uj7+qNib2n2lAX4+zM41kYxayTpPrT7vonOsLPRJZCBauUl8leXovxCVdaFFUsNrowQ7NyA2MQlG
NpH2i6RV2vcxqKSi1hTi48ay1hMSGSNp7Yypkj5fjBv/3TT3G+ooFDPZz9QM+QqGHTGXHwL7yUWy
+4E6gdmMlRyAlA51ptoqwNZvxRKRrCYDYTshbmbzd/6wBGLnHpbn2fEffNebHqXPCHaR1DpnF7f5
UwsXbCQ1LiIzz1HX8Vt6hXXTt70gLjv9jvEbXitPwa+93ESZXGnHXHD2b93IPtTmKjoBxw338j/0
F8Mb4xDeSqNtbTRpfmoqRvO+/Pte4b2e63FUANaqccNhLQAJ1GYgK1Ipa5Z+T9hgCtLNiqx/nprz
3ATcOCdTbQs64b1vqDrfpHOReF1v9Fdtt96jEgdcwzVzTcYLsGa/B19Dg8K2rHxyh4a9ZaGWwuTb
uc7w3/EFzqjpaOS//AWSRm564Qqz/FaBDQT8k6IGGrpYGUvjR1sPzGgkBSeXRRr4IbTl5dw60TRn
8Vm7Ur1XJIwbmUHqi5cLCBbIAACRM+OsM3mvz497LTjWWq/P+1h4Mhj+IA6Bs10YebrBjlPwWnOX
rA7mQS5D7CF+Fx7Ru3nHl3z1MFo7c/SigN+xAPxHrycVcRYzC/tDp4nN4//zxWmxVcsXvszY2zhV
+gTrE59l1/7SvAE4Xq+4LycZ1EdvjSL0xicEvhy037X3cUJgDgDzORcxfdSJAasEDtIEZizI2K2w
AXpQhYZdv2xDLtx0KxoO3Q/ICOz7wGOUr9y6zxJe6+LGwoqbfLsxXFRMbUO/IGlHdkJ2ArVEzYDJ
2OjVil1wkJE5raWHsJvgHXP9egogZK/S6MGBk5MYqMZ8ieV9lqOcYghZQ2sWutIrsIeBKf3/fdtn
i+6VnOEdx7CoeC0j+IVD7lQEcI5lnFE4dLBTK/MvGxbpzJzBZKMqn42AGNWG8UhphJnvOLEiEZbS
RuzZFWLOJ0ZEN70YP41N+HLO1ZXS9KLq3+MPcYNfpUz+QIaK1qc5Gn+QzeGfwH4coxDozSv3G3S7
pJSWMffwQrbhp7iSc4ZTpTdqDON1WijQTvpfgc3jCE32QYxxb155Sy/fmmbf5Zc1cSKuy/UunUEl
K/0gFrahgn7NvPF43/T6sJoiYDs3Di/1wP2PbR7Q1mlT3qRBWMH670VEMDBpdGzuQLSAnOv3LNf6
80WEToKlSmlNx9T0nI0jp9qHyRprjOfeMHaqJm1BAvdSpqeybMWwdt5RHP731Z/Su/BFcWcjk4lg
8dSrK3Vmw76SVP0xSzmB4mz2wdGAyHIQYDrMklEjw8enOzQWMMj+mhj6b8LzQ2iKbzoVsEKFahWk
rJivpxAgxe3ubERzvLgGchCU2Y7+wgk87vYW1noprriZ6IQwDT11Bo/d+8Gec2h3fOV05TYqPb5v
Swen70zu+wT87iCVqbLZUanDuJuJZsDJEUCAhIo8JCOXcXhYr7VG2Z6XAT6mcJhJO09OlTSzlw+r
WIpfAD/LcA5Ptk2C2Sl7MQn0pz2eFOIZFjB7cEo7sHnP/tOOZmcmqFyPEYO4MS13dMGRjFzcj5Lb
HYSJYY3e+9L54MeSy5yNzQabQl+It3BoyatdOpdSvNj6s3NwF1MIMTTTavHcAHLMfcEdubFbiGJ3
Glb3ofhplf8alBCianMQ6dj9BEtjsDRPyivJXN2EQ7E04mZ9WJ2gcP9xI2Ho7ydyVx9DZsz/52rt
LLw81YVFl2nWfA3FLUl55mN4tyPxsgKGDK6ERxVsDUrcLEp/2O7W5Zqs88jsO3spNYLIQ3L0ree7
WUDYovObMEflQoSBMGQISPY7KEyoZTMnp+unDUBPfXU8fdxEtcbOMBv4EJED32ZPjnTVaNVKNeys
GNkyAssAtWx9pa8c0fb3nQksPpRQFZP/vUlNKP053AWAOXETdnHDkfZ/K9MWJ6yypYgUv2rdHfKu
YRw3kuwHONhrSPjVh413X07XWLE7cJYPQuwCHJ2jMuGSziYCtHKZCxkk2gjny73U2EJzezyNLNKy
qgOOP88P5bfXbTK5xpFI/ppJB3x2Njk/zJhLMTQixjT+iMp4212miFfz0/fE4KSXnZ5E4QNqu7Xw
wUgl7LbbZDS0CkjWKLcu2kA85QPcCYm0Nacj+WIwmxV10ygsznwWlnCb5YvkyOBFX6TBOKkiIHLZ
WbyDj77OifmwIkLUnCVcaoeZi194M3/WhTfTCsn+t7dLlGBoE6Y3xgH4H/dIMeEr5oCwhAQO0ffX
v6/F3m/LTfyJsUZsqfC59lfA3HUZQQPJFxz6hdmj1PkejKBS1ZIPkoIz3uhpNsmkZT+DGFkcmi2y
0o1S2wyt6nEzj0qnP2vcmNVoEvvGbrwCrAd+WZCdFyf6SlAAXAUdJiH/pKxCfVc6u1AjFKHcqBBd
SKxQcYDssoycKnKM2DeoTXOSTP8gpClOtO+N4GDNNS85CkUU937zSFYBPxvpRUfMZp3z18xSmUUo
+NxY8N+4YJ05cxVdzMoesiHxQ7Kh7BUYYT4OtlU31GlSdW7L5NBo9Y76Z2fYTYrb/1S9EQhsKJts
Ao3PHvPF9gVBjBM2KIPAwCWpnAo+rib6Mj3KSUXARHyAqb9D6I3Q+9NR9nUer/7d6vSbu6qBajGq
KgF7Qg1hVFT1duTyFxKzUkazIjtE4oYYq/ms2Zjur7+yJFVRypdAnjCt9+uAkerDuwEBV63eFHHq
Vsl/SWyCxXe1jYb4w4NwwMfpR4Np8E9AUqUJq1u2WEEi0WAx8P18CEfwrIKWs4Y/iAiHokh0nO6e
zpK2cxJBxUYvEBMCCB/BbVhfXkDXwsufZ+zNtlBx2alzfAvHETMtRxsEGz5xYYNDfLDVDYuK/nup
VxCMGmqWjGmXtUxxqMos5HdZab2WOzwXiapYlYw9l88C7aR+klUOsJycx7ImFcScjHz52bEASWCD
nQxR3iMeVZUq9iJjecHfiAen1qy3SvL6GggOxmLY5l3qrsFuhK8RHj4DYSWs/1jmy8Btj7LqNJMH
qx1PhlZukpmaZTAzKS5aXJP12qp9SXAbFAP8tXWuNDkEvHjAV057wNHUs3YZrMQGoLJbGfr6Xijo
XrziiFsOxm2ygzb5WvEPQYQDcuvmf7Xh/Nt0AFO1fJyI+x3CGYA3yUMCHC5/lETT5t/0wpfwFdoI
VaMARf9spllPzfj6dcPaxZ48d6/WIYbljyj0d9hXgqzEnYLmDuJqFek6JnXMi7Ah3AIHFnk14V/Q
VVecO0tdHKu8/y23LWqJXYUtjyEEZ1dTrlb9ggMLtFP8g06k0m91IVrViE++oEQoB07+4mgHmH2j
p/JOon63SCzaNvxZOnhztE8tzfcUSYvq3BBG2HXZDJgO5a/mXN0xT59uTDa6G+kJLopB6nwR6ROl
9ljklEJ2zNlWMo3MYFiJcdI3kitc8mswh5TYvvY988IbqAy2q7Mxt0duaWUizWUF1uH8YYClSruD
ubq3AVR0LrR7gnzLp5uS8lkNHDsI2y610oGTDlq1OtH2eeoD5lXXnwsTISTLf9MGJ9eSLA+1+aGI
x/6GxnVrhU+Ht3JgIuGh10r48bbFBeAjuIr4hDiKa0lvHxWNfy4sfOieIEZtAJIDFiX3kESM/I4h
BGBq5kzBwVBwnYxSkTiMF7vAU1E0Yp6xrCgu+i02PLdkNg2WLjLVDV7jMlnnLn5lvf1iGIZcj8M2
fUDhoJ3FpkJ2AzuaHF8xP7fgng8K28HLXPjl+17Z8NIJmU62qycCSy2vvJLD0uRf3J9G6whAPiHC
f/PwaSWmYtAxn/kaAOrQfH2nvDrP0FVl7xDq11QIgIGl4zxWkwioMpC2CjlVifk7+c0adb2Rf1eW
wusZnvUOb1JlLiutBwMmfm4qSzD7wMTIetT2MeYAZGNXtLJtzO+E6xXjHlXWoboEH4dtrQuSwPuh
klFo6Wv7ADgOGw8/bJr4FB6ZPuy4AFKa8rYBboQswi6zHKmwXbuwQ5heko1wjRURTetorwaVtG9R
o5pDqIwA2YWJBYTt7qeAZ1Z7V6TRJo8g3FZI0N33aP3IaJD81lZHWnBzJ8hOLjztr0AV4xF9KbWZ
3C4xqus5nW0S9hlQAiOc/sSMeP4hL+/2BLa+AVACk4Riph93cRxuYZdj//Ay7z8PzUe+pKBsKl/V
dIK6rsSQ3x7V7kVj4Mcf9PcNdBPbQKM6KurVN6mDaDNLB8Cn/g2J0TNo3zPIme1gocpYR/1deBdt
kxMYzLDOZjxjxI0EmOT3kYvKrTDlOTyTIiUCjhIHPYEi15F0KDFP5Y/qbA9x70CyGj9DCvFebDC3
/+cuJE8qSWemm2ByjYyLzLKNRcH4Vs5+p6Nbb5bqy0vWmsfl9RtDfgjWOwrJtOzXo1bFJoAMrAWC
+K3zhWJ43dd4rkPlRBNtS9LRBplY+olDMnNSY2GyKqAxdSHgQ5aaJih+8E3k+UXdLFEk5YTfL2gA
lYZKsOAlzFw6hJH8dGuBgigoNLQJLHOdJM0rZ8Rw2hs35N+vpGUPb6S/Jg93TjXXjWWA4mMecqRx
JE+ewsZU6T8wIGl21b3nc+36kxjKVzGQ6XQAzZHmpWjmQKDPHQm+83v3tJ0EVhn/FmyunQjTmVKg
qBJG0dAy1lJ+o95bGvrLLzOZlWaOZ+kiNeXU6nL8CFzPUW3QgF6xYozcZFH6ojcHQJsFSDoV5dHg
CiBtk8KA7iGZ3Y0txfoe8fvxskrFlJ78SDWVYicF6A+Du5dMFYA9xXVotkcbRz+qdH5iOLEkXVTx
4PKdj1DpNcMjaZl0oQZDe9SPLtYt5FIduGvR+vmXJos4PqNwmYzH2jbABnESXabeNp/f6w7C0hhl
IYi6Rrdzb9AtjMMNulgPvNurQ4yVOggbGAdEJyOYMNLitHbv0MQJRSriyZ0tQ/vePY2dKtJkh+hZ
70FFHEeBDf/gMcIf/Tdx2mNsuRCOc+5Pv8ycs45MhNJfW4mrAMbDVGI7r6ZvGfjfamXvp3JxpGrR
dJyIAQ2MmwD3O9tiCHJwad0ps6qoBiXrGbgHWrPfwo8vKnuKbCka8XhuBmCk1TiYmvcJxstGXg0i
VMF3u55Fff9KBvEKYP5vTKF/EDIKf58DhDDwzZmtg9y/taWrVKu0umlcJVRIKTHmrSudl7PROwEz
bP4/7vNMUmAlAF2Gz9Cy5BO6Eql3K3DMek0lSQVR7y+16xf4GXLM0UM1daHVR2VeeQ22Z1eE5M5e
vPMrx/WoIxbZVbtOVzqq0AxHX0qfVpp9o3ja+OTePlYXae8ewlTPqF8q7amEOc71BFXApW1sqHvR
wzLxvdI0w9D9C45i/W7cYP4dK5R5ssJXYUdbc658dNA7f7Kk+G7pChhYh5yKG3kjAHlw7oL+icdl
GttLpIQ1heYRY9Eye2BOFY9kwnFgqY1iNFrqDJMgv4lSRmNAIpUZl0iWo0ra/+rwoxkFa25Zt5dp
/H5Lfh3OkidJEyP7v7g84TN3TcZQWN++2QMJlY8B1qLJ3JqfJ9kK4p7ER9eRn+yK5A7qR8KNaoY4
boga69F5d0NFR8zsCSngWPvcArSTZTk845SueRAmaYUE9KFdUPnUMYeNRjXCP3OvNhLaLZqFaK0z
XAhxVpzJnI3pR94VoUcPISXTKNLgqltwLx1AbNnhAm/OzAnjcX6z/RyKx5c7WiEKk62ZN3tL6Rfy
Ei0+Rbsd7n2xUh6+n614NiizSret5ipKFIeZ3xlPKxtgsiRd5o7WYbAgWv2Z0kfqxgdNBM0aHroD
Zy6DqMiu424ab1nHu1L4YM4MiDfIK8627J0i+4ufu0jOpHatZc2VrYaaDkPkUc7bVXAGg4MbuddD
aO+tTs10iWo7JgSZE754598D7EJWuVEgUz8XFdRKwINokLQI0WP0zZ8A/Bm0JsoMhTOBmMCxGVFh
+/L5uscEuRPbfdkY1RxQYo8Y0cQnXmad+uVYB6G+UGwwcYL6M1vdN6o4mI9lCMbKQsMZp8jEbEm3
novkGJ+sjQRVxKDL+lyzVVc5CN/g3c0utcG8nFv6vsgcL6TeoeOYM7Y3Tca+EJsRs1/WZtAynpTx
uFqa2zlnuOsyvsEptA6pVw0cc7fxrTWHsgAaENj/osvni85pQYuhIJ2TZ6e/Okr2dios9i2PlVFK
VX0Ak+/MdTnZmHXUImL5V5ZL5XvIX2+FUIt9DnG6182/7qHfA5QFADq3nKi+m56R0XXabkSO3Px2
9MnkhJLqqEWbZIJLmS9H8k64Pr4SL03z2GG/ObSoQHC507bqWX1VUOX+XZrKW+Bo3W5lCaMVTmMR
FAyt90OApYGmuB6szKGN6Wyef4HseqUBVowyJ33ooMOMW1ipXEA8X+c0PKUB7RpeFhXyQsquoBy+
D2LmOKc/eN2Buz9GNnMlr5G/s+7tpPtA1wD9aZapCS5B/tCBNGHc6KIU6orjVoKf7yZ4vR9K21pv
Z2x9aWxJEVlcEOKvpdrskN/SrDxZrItBPh1Kkm+sTiymyLdjQspxnzXT7nR1awx1ZEHcBlmORgbD
sdpqOJ6xiQVxNEN4+JM0uhAzUzNcdZZzmyL1KOWTqj6qjEalKzqGevhDtsqxI9J7us/Q9YfKo2lM
Z1swWD2WHWzDKgoN1gwGVHS2/V4mHyYVg0xfBxdzTjc34NacGICOi/yhDME0KngaizQ4Xuu/KCp8
AJFvSNZxPUBaM//IdPcdZVor/wLbD2wa8SZMrV9ixeBq2pT0246fSF/lDQEmm8Ef1Slr5BFMJUKI
KJyrwi7l1m4P5RS5aTy9xXHXgIaW7bxIwFiYWeGmdKukAl7moNDis/204Hdaj2R76+RXjS/T+QP6
DPpEWYqcc0uVAAYVqcnuM8MqvGQstGgaayow2YZu7U5DPG8HAeeNih+SL47ZOFc4yLq1M/FsT8d/
ap/4HqIE+Lbuc2mUBCheyrbkopZ1AucAOP0sb5sOchkrTMtTSaO4eXxXvBMp5LyFYqTO6vjDvHds
WVUcOtoecHHhVIUBpJnnwXKGNuqTqeFFLinSMJNxRYEd2UUBI/Q6+/NxdObXz26G2gMzcP4E+d9j
WmD5VeViyLA+H5Povrp3meeu/tQecqjTsBcOZareMXE70cfSYRMrBiNG6jPWv3QKiuEfvGwWAg2E
J0Lae9PrCS8wVqnlQxOAgNDNU0pYlc9otIQlAdjRE9/ppq/x4rF05eQ4vUoLGPYgfoEUgE7xC9tZ
+tEWdTUQlLKnasDmXVGMPUH7Bj4ihnFUK/7subz8c4oy1n7lF2Jy4MQzFPk/0A2wPQu7aiQvBO3e
KkVC2ka3p8e2KdEWBpUIt4HsS+22u8CpljJQKxVth70mz5Gycko9k4x2cnn1LmxDPDGzLIAnCKD8
Ob36rEvQnplmUFRz5v3/nrFAO7tSo2QylpHfOieAB0ZSCMA0YB7V8s3/3gBe0rEknYeru23f9/0J
cYSttkj6odHeFnlIuK90nvRXv5my6KMMHmCSXHLxB5HhouyM/c+nXXFynOHLXNrGdFAByvttUeZo
PZ2pF3HiFeLORF/Rpg7MTEgKMEYlwDGSWNqIWeH/KbGkas1ieKMylQPW8MXAcx2WF2KUvQoudrID
K+V8o/11F2aEGnY10WPQiuVyjToZHPDtB5xJQ8vgwucx4UUMURMGPtO5ZLhIPgdECrz4AimXyzoB
ct72HYtOWhpsTiDmzazjdG5bfIm/OURWo316GV4iQbrI1wmJonoJ6x6sYoXVPXDoLIxgJfk2a0to
SwZweHXEqKgljl3DpFp7p4BYptxRuGOhUYgMZJphHM+geOQLDllDXSsfTELj+e9uZNHKxI+tG3PF
bT3QRFsOcP3vLVGMXoX2k9eCPtETh5HEezbXFguAZ/n6qq1uuc1F2jpLiFyej3d3eV1x5fYP1yz1
Zm+YTDMGPsjePDTyJ9+YOYBz5+PvlEhJT4NmYxNxpDRwjXDT2b59FxNpJyCO4uXO8MrlGJWVD5u0
CzAuXIb5PUvb0rw/jfy7TjPdpGPKp0RcqddD0nV6Xlkdp/wNhpVzcs9SsNLzB58EFDhoLu2IIa8z
+xHuAYpCjVGKkWIkNeMaC/jWgqdk8wCitgF2dEGusVFJJoVpREVkqQgCgBw3kFOxGBr3esQBeVKP
EAHbE6wFJ5MDzflBke8JQNb80DJalay5lv6OMxfLu+Btz3EJ0Aipeg4TD2y+zMbwcxjNHFAfK3Tr
6aNt+lWlKztzzWqEDQbBJY7B52d6GoGpHjIp3Iu9z2SurkS3XPZVNGvzZfnpk7/2AHOXxBXwXAtb
7lSNuqGJkUm5HHIoI64+URFye5sjExE0Vf3vc7qI3AX3q0VOmocPctwjkWegwfsBTYmUIdw84bRB
eaVdo9fNndQUF2dkNqxmZEvVi3qlQp6A07AVklEpiIKArfo7v7K+JnUAhWxP+1HxioCrbg+qTIdz
UwQYlRsoZtA8vcM4/eT5ATjlPpCtBab9KtPosVNQ/jawm8YcX7gnzIuCIkW/OWRUO1yRN4YMEieI
KQsvoLIwdtVqtrDj4P01F0EQdSrsRWnG5NUQNDo2FtHjlv5wg3d+4Zqs5nbbM6yp/xZr5OjtCHrC
BbcQuEj8Eb8k5rA2Lria7X2Oqk3uyjksbMuiOPHY1ZTr4PEuImC9B/M/uiP8tWpm8zl/R4enncH3
cWN/J04XkCuJZWYsDqrhSu0sa3Kt9GWwwZjLmu85oy1SWBSHoVEHg91sew+XcZ2ptASivEiPaeic
pVVgvuGUP4PVqihcuJm9vwMDiaxLp4DGof2Qecup5TB2mfAHU+x9pK3HYX39HKGKIMsIk2yA1iwl
6H7haYAV1xF6K2uTQyK07+46MRc9+4gv0+8Eu65bAmzAdmoZVEHwBTasYYfF27o9GXZUWlo7ZumC
60JBNufdFlAMJJH78F9acQcMXIJUk2duqmMJAbUmOvJy5ff76I7zSM0PYAJG/R/5FiWZH8PVI6TZ
ha5Tui0SdFT05jrzuevIgRCNqlaEQkJxc7hcdXxNt4/tK4H/vUXkGz8xEOQAC8ZkZhe0gmOv4Rhh
1jMF9tdEhFupDtgO+O2fE7tVi3wAwQcvUZxnvyQHdjqFaJTFmkeHwnsm+QV3dRuY9BKyh81c0ifJ
lQiWdN3aIcJ5gZm3vzjL2o1RuO9n/1mrOsK7ejqxLLefXRDdvPRP5grTsXFBunkqoV8AHqAuqhbl
Ucv9GNhLVNRjkUSQUdBJ4nT8mj6unZN15zWDLo28LcgZ7+Uiy8L2Y4BGkRdRAlXRda8pS8J2nYWz
nSJyv9XEPFvlrrwLNI3cMmksKtsreAjT06b0LsCBwZD2IL8rYM6muCf6Or+dsE9fJcx89QDmRNLZ
ZPyltIqrLuqjfg9vF6MXn5wNRpIbqUB2FusQvCOiC17JJDPAqg2fslLNrvOxgP/ImHkWc0w1zgio
g9exXtG3qzeUPuOhzXiGJttUfT120tFlQFOQ+4RHcHxyIZ8td5sdl+xYQUxxN/7a913tHPt9x7aB
aJLKPiTaFlUE/i6lnwUgR5KnQF72/tpE6v8DJGgVf12mSqHINqlCpHpc6rW6u14ycFv0Hd/CNDGo
kr2WBWK/SfOday2UijMEInSkogikocmtt6q1iBt3nITxdY3yqpdpJ2ny6ZiCaMPXZyWaTr0i6jjt
UYP6c+mri8Odt/0yjeLG/vJtCgkQAHNz1Dtxzw0FST1TGSEaY976hSwSRVSpZ75MvJaKDvvXD7+Y
2HFsyB80UFMKKsXoNQ21ifbHpA78ov4mxN6LmVpZY5kJN5m0qb4hZeDNA9TFou7eZu6Z2e2re69y
9XiJW/VL1u258ItVpYFVxLwilKA5jI8qrIwNINWnS8/xVLJFneoFzj6ImyY2A2p1wtSJT1lwVjSe
jWHoDUk6oKvX+LAb44T20+YQ6JgwpyF8av0/KDbSa/u31KRXT6C8yCyI15Al+nfEMUTxCieA3IjQ
9l0S7fAW2EJQvHSvn65ixeRculCJZXW7mpQa5IrcYkjn+GsaMhY9K8FwxMl7/343fYxpnUtW9TU5
uCltYSgJKJFCTAAsmWHiNcSZ7ZQwEUV4ipQNW7fERme9g2qSg94q4HUAAFN8OQVlcOFhDronIhT+
wgxQTROUqSClRQGgjprFtvR3i24DiVryrtDgyDNg/Hus/syK11erSYj9Xuf3HxDhFdbhZIKldMLn
LQz4V6cgys26o7MqYtpDOsdieGv/ePcNJ3cLmY1r/K3e+sGI345CsoqrmM2X54nLTxQx9D0ZXwub
CWY8iqmC6Y64BwX6TZ9gfRXvi7aRm6y9yJ1O+2uhmbMSKg5Am+/pGa7r4FT12+XO0RSU4p9BGHC3
pQaHJ7bGhPGfa0WIjsqBwzZuiyvBFbtT0pawJgdcjMkTovA56d6p2PBAFa1Ele1/PqhohrQ9X4w/
exLpTKQjwW3/9MYTohpLGFFHrkot/4VY+xmKghq8eXAoXBJdsSz9lPynGnFhZdEkCDwzU5DZxHLn
RezqdvHRHMdt6V/27kYc+4s41x/60nvlTtuq9GDUqShvBY6OON+VGF31UlpwbhrX26T4UB856Swa
ikiCN2sFp+x9yoOmxI56fQnZvVecULG0cS6H0sauoVHT0eJyokZjva5Ye7/nLWIUnGMOBugsiMHv
Xds5mnO1Kb9eq5wx/h2kgASVexxXP1urQjSp4uF37EN77GvDF1M6QLvCR9WBAlY+JFA+WHehya6H
kTTZm4PI6IjQF4GJFQbPKyU2ItsMRk/VgDaJBMUyqW5YHC65fasg9oxwxdnoKUURKy77/fwnJGjS
cSgs1Isg/X9d6UJ3toulQMEKJ/culFQJNlK+tWo4MZwh1FWRn0cpQ2XaqRzlYkd0sZzluovfF2mJ
rlCYNqbHUIi4fa5+vgzEDB2JbrrRY9iUh0ZUZSVxStd2dy0U2/kaT5XtCiuxqKTc4SbMaTSTulp7
kXgxaxMDGetdJdu8GoZB2NMeubsomeC0h6wMsnqt1Qz8B8fEHiCnbmh+bkjWAxQGzx0EqJ/IugdV
+jIW0ksw0+qFr8XpZ/U1tACrqlxCw0+aYDsRbHvBn0ieLy+FC+NBAjhnAo0Ta/Gj8aGLnxTmyvfy
hrwNPoYSm1riAzD/SR9ijwx70i+BzBh+WQUbxMPUDC/3CMcXn56UTah3f76DZWr2Qf+m2VeJtFDs
fDN+XoXiI4U75NjP2lXJ6SHrJLtuuMiLqt/uBGFHXbiPmBzWD7YOop4+Ts9RvlsGqiMUuUCjoWoo
bf4zYuHE56wMmL+WT/6q54EVZLfXwRSSqNi94PYI573lXSJexL9zLQhVAcTwNuXfok28UaW/rw8u
OnNMbq5mjscY/IlnFNYbVUlSjGvuGlcXsgvzRu4PLrzVZv10ODc+q/ZlXIeR2cXliev8ELSjYG4V
yLwfBf+DVEk4g1X4ODpSfMYT/s2YdRnTgROFQRsB4S2csD3eVhzxn7rOB+zxD9QqzNF7z+DLklrV
rtJf0mMl6eMafX2XByacHkqwUuKDMIQocsmF2uKDwLH2fJAZ36me+G9bB7GoKM7GRRYWTVjTc+qk
Yv0rAIXVY+RUnlIzwDy8wxg/J1GOzJvCRXiSC8Y+bN8IFEx4vAy0ESWlC3zx5CGLuw5Glo5vFoUv
s6Epn/ngNR9pdjx2WCHh8l2fiqB9tfzMGnNjBNNCSZnkTlJmPvyxeNKNsm08rrmFQ9FNScZqhW9v
bVjFnlQE9nWaXfMq/05nX9VqL0ad4Dil+U8VfKaz9m+1tqxUxB3nOhkEcEpjUxT2NoG5WzBXmwgC
H346MNQKVfHzVt+3G6QJ1r2hPhiImcMTKdCqGAK2jEF8AmJ4PMDR8dP4qXApuKCjUBqcX41Z2Vwq
wC4CtAKS8LiIW63LEhG/F7u/DD6SPWvr9b0YaOEL0QfX/93ZDrTvyM7EwrjDuDu7WB9ZsGifuaQi
sxGYRkkn0KKZAbySWwDjKQn6HPcb0rWPlJdtjLUUXvr5R6BP5vXCjqulXO/zKQvg0qBKnH2UjSvt
H+qdNIHkn7sK1EMkfY+46YwTCvSIA1cPmC4NhMi+jz8Wdv86wfLLG2aqTIfuLxTd8V4ZugJN1twP
qf/Q24Am90BXXBram0+HHvtvWM2lf7b8GseIgbrHSlRUa+BCI4qdDkGScoD3xZCshULSUhlEzWom
t5iPHC4+Lgre8kNygY8FI4JttBPhdvuwmCOK9xZkNOtPeTg8fiJkim4Fm1QvfUYvyr61D37b+pyk
s912i1ggah5rpI2EAuhZW/MSWU/PsRpFAWPBvnQjwVaHxX/8STmOtPiKsba2OmfCRoBkT5658oVx
A1JXIUTllSxf6Ft+OHObXUxuw/K6jZw+NqGCs2flf43hlFynBBMJjYd5PlLmD2tGBWdAK1b9vihr
NRUJGnExsJAkij8B7OKdQBoGO5WaeZwfvJzNaxIO2fBKTRqD4+BP7PmI5EAd+wjyl7XYRKR9LH3F
vUXgG6c8vASFD0AYXBx4ndpUkPn9SFrc5TCYekwEKZ7PnWy46MaIWvUbklOWG5fSmYkrZmFUCS8v
GN94waHFr+C8QDXxvwAxsn2Iljwohnj1+F7706X9EbD07nB2bFPj5poH8t8dVeR0pKV9SJUcsrd3
LUuXWqRnPlRNiQcTg773pdkbMHOHGU6esjhLtHJFmyNc7IA5kVPPq7xJsofkdYjRvQbsKDVWyyl5
lY0rtKCMvboW9yYdErB2mwzc8azBNpAO/eJmiW+BhgBv40YYrJ1wRZ4W5MgIS25TqRL8xpLLsXwE
ZNRuZW8n5YslPY1bNPUqKoQZfS+rmgLuh8iDgqynm9/6xSifRIQisGTfvjSeCR9B6Z+EJmMXG6tj
Mizrb8NV47P6Qkr4ypvrfohKiRSAPbO1qfAZ/kFjXz/zIzaw60Pk8jobI48ubEFhlV6d1BowTUVB
DQwejG6k2RqgOdzGEuamMny8GyvfuY3BkMTzJjn6PF79Pz6tf5GiOj5EwJ9yOCQ+LFK7RFZaA2Sm
kjkzP5QxoUzY0LFDomcmf00VoekUV3cYXM6DdQoNidJsO4AgZMwqkR9M17OkuFdH0NqAcgMC1Slo
WTiens8MDOsTEe9mq0TLXGDux8556u63IByv5lk8TjS5ZKp6cZ0Z8NG8xjvGNKMPyVYXw8rUIUpT
VdyRQdY7XzqBv8rfvtubE5sMUJePgantu8IKbhrmne/9zKvdlc5iiF9m4T8vEBFzrabLJjEn5SwV
XLRZcEG7dSkWzApl/KM9WGIPapsEvBwbsefsxrDN48wB/WG4vgA7tXsF3vK52xZTm2o262DiYB26
o9M3a1hiYxlWeU3cVnBy+e4chZ8dYbwanSEc35czIC8rCuZm0++12PPngFjuLlpNC2S/uPvFU7ph
ViWComR9EFsmXlbOew5J7uywCZMtImpdRM0RYO59G2Sa/FXdDPJjgSCSDqhGzSJnAOP4VQnLRdFP
1m42SLHYD3G06ANLe/MA8ZZ2UXqFVKKDe//i9yjLignD1C8VLHZlua8ltQCyuviefequsFjUcUjQ
sKKjVwH64qPo3zSBVfSB6VhKoxmX0g0LhPxA6e7sKchfk/zJEF0pbP1G2DlKu3Bw42OjbCm+GEEJ
yFwCb089gegalASI8oG8vCMIef9IVTEfe2H3YbvMNge19JYQqUReHR/MKBv9B1x+CQ8vI0nQJouW
gDb0XZqE/AGTsRksmLRgmyfIqoQ1c7lUEx4ROlPX7meJUvF6FgcOf20AzUu/0R9pUMv9JEmUHlQg
nkGUj3OvacP1pVwjvsroWzpR/5DWCmC7rRUnsuLoFuC4Mz0KJ5/jFRYGmKEa+kr/sPDYi5wG21mU
+43wWo/DFTjhRASStxPuzR3frEuukfT/Ezlsy50uLVQ4D2Z1r+LcnXuL8FexSmpiDnJ2deL+GvP8
4yiVCvxcD77TrhB3HiF1W50OsqWw4wfYFqtTN0s4QAGIW5PXFVRiD+qSm4n58fJE35+BDFW2QmQe
OXI06L9d1L3iBJU2nP7yjx67RLNjLb4tuEMyPls3P5gupyaAWApvas0iT35SL/rNmSR/RvVRUXDR
tVAHmJqUWqJ++Nd+EavABV2O6rAAGPv7vySxUWc/cjXT2Uvvct2mqD8FHYoKSgUW89IoO+zkG3GO
kQIR4ld4St7E0mJdfq3KK9e7AhvHD656YfLWqVei/YlP4p9uZOFcDPCBtkhhSAK6nvelI8nAO8mC
OsKw0wG9nT9sAiAeGUrOez7XjCUK8GDllRLRJLnaiUeciWsU9QUtyTVJtTxXNZ2EnNgYHaksu2PG
YZcDM7huQ31LswGKDLuFWEpftpfw0tRrgRDkc0PAhgEuQoFOSJHZUD/zIfJxBteABEZ60lsvgIih
2aEK3ZwoKToeuEj+HdUlmntcE0pH68p7kvinWQqUcwlg6YAnlCq3x2pg+AJ7227n+csu4U8cU7TC
2H5GacMsfy0tBKzwNjn8Oc3pf1FxKGLaelFJjszJYwGT9ka3GzOwzkofgrFCWozwtgUUbrJJO5qm
Db294d5TtuVfYEGdAm1FGAiKOjXLiJNDsceWrY6O5cZS8ZBQr0YxC3vziQU1HrGoX2hEdeqcquYj
mVMkNHB8RxNZURC1WHPUO8Fv/uaUI2YtiPkHh0clo0Hh5awI4MmKrfNhQFCiQgtLiU7KwVnVhqz+
bszaYiOVFn3xCu6gJ7a3zb89zzl6o9DYuWXJK4fCm35BxjxQrwHx6cO/hiNn2+WjiBtiCG87S2mm
gNSifalGuQ8Tx4gF2oGOi6I0FFdDKGDAit8pY6SkIePWldiJdQRO2cr+Rff7zin6i1eb7zstHxY1
bQym5YOdtohN02RGLLHo4LUVTZIlZOhgmo7qWG3HujQXOaf8GZVRsvvIpZZUhn8juUHsdXurH/3u
tF5O3FtZi6l+vly+tjOLcKYys60/KoA6JmXsVBMxKiM7QN5RGNUC1tKjeUh0KyL7QIeqN58GypfO
dUinPT6V9Ga1s04rlAwge6w7JSweKUhf6A9Brr5Ht5vtXzB3YSuwNPAGw4YR7MLxzivAd1Dm1qZB
X4pTpXH8BM2jjKz36skVZ4WyBLAWlVGFCQziuTy8g5DNDF43o8Hx0Y5xQ1nXpdZsS4yLoC3i2WV+
4wG71h9aC3XnkAWngjDQ2t6ahMcHDaedQOFVpZNzIDZCNUCDxiMPvKrqIZ03qIDS8IS6iDrNajAy
nHBgA7hJg03bM6Mv+HTs9sLO1sArtOtj5TKjw+7QZuMtDLI1p5SNcgZjpam/R3aP6+heU/DUZpCo
F80necaxGcZefaCF36EsvgEC6iETGIG/ZmXM2a/A9lQWjEOFudeJLWPuXwa9RlpSlZ3LcjxOilHh
cASRvjrtI9N1pS9nNWxAU03V+Hl1A2W8WjXB79jHGH0NRw7l6uCGOmKupRFqWd+dSOafr/n89Y60
zZS4W29UBzvZbrwcLqjhyOQGEMgP70+8WDpNxeRrTMVrVHa95rLnhn6fQikPGqAlTPsWVyqOJrV6
oGdTduj+gK/UpP/ov5yb1N9JKlA2l5XJCGAggHH8OfJZiISQO90o4A7Gl7Ifpz5lVJNavbVkaq5w
VJTPU4lDcxTdcxAntzIZ2k7IUYmKCKzbUbTe+DmfjoQxg/unAG2wn8dN3TWE/yrjP37h9KDNEQ9V
qzswRro2IFsIfV7IocH5Vq426+2kgigDcTx1P7aGWj6p/3E6rJydH9UFFAo+hH0uqU9uTIW+nKrV
46zJi/HsE7y/Fg9H6dzv2PTSD8nG4MgQaxAvoyr6XelLFwkU3HTVkNOy4ojqA9xX1v1rfmTyAss1
pRxgKQPOpXeffTZ0L4T7An1xB7Wr8rU7DQUzS1GbUj+gOsmMllfgzNGLUQaEj7g7mYJ3CmKhSo9j
fclYkCxKbAu4tRV9UXzAMLcEW/gPwh75Fl5QLAqnf0RkTR1ugBbcfPOMzHZ0sxU9E4KNRXoSVDbk
9uFJvxvqQ4+5fqJhmEIibTI5E9e3NxLC2Jlq05oRrQqE4/YKoAx/kJu3zxH74kNxwUf9+6jomXBp
4bbM1yrU+iqFBLmLm3Tvii2pTAp1JXTk5KjH6kNp0Nw/BWLZlKDpPVrdmNhR/Kk7TVXjaZr0H5y/
ATYtP5QkuVkmWRecdvDgrF4f2ouLH/8ppTlsIy8Vqi1qqMUea/dPImY//r5Cw1DWz9vDTrGuDvws
Y7x9Pxp/fgTdzs8Q0N2r22Bh1ABGVud4/mXkQ8DmfJ3Kf5OPSgk2cMxRA29d4D1MHYw9py/gXgVL
Da3d1oOVU0F78ajMHYdyKOQU1nRqwx/8LPEvtZZkC+W6ukMzC2VXwsB60Sc2I37h7HEeldT8YaGj
Neu8xakHiA2KkEQDusSrfqmWcM9EnqcYj7UEL0ddOFT0PohoLa3LZ0AGFFUNFAIaQWxMDEWjVdwD
aXQ11uLgmH7J9aiL7zSuNuUjDplJYoiZ7WrNPhY9dNUuTyaD/u+f3h3LafWbVKoQ1SYuFWxk9ZB7
IGjjo05k9adc0aeeY4v70uPr9WkK2fWhWshomi++pU0fhccpQl9TQDZ+O8BFSwhKHtV4w2rDmTia
6qpQMZ54GZh66QTOV/q/JCP1Ga3tbDHeQAgIH+KklGYWOMZqeDBaUNa3ohvGPUwUXXZKJY8KnBQM
CrmNZMtbM/5PkGSECstxe+b1HOc76Ev8uEtbDB2E+dC98zBwNyCJZls/2gqSfgWV0Y3ikddHTFDv
cOv2yhj05/5BLQCqvf94A7OI3cOGBvt2o5gzVhSYCG7grI4GrGzYhn0QMNXufM7f8I3jm66AbOHU
A+6ObaZQTgStoFl9ydVP9zlBSGhc+efvkvKJBX8V30fvmbJwFEvhYGB3QYjXDZZD3ENPh9+DI55I
7eC9WaN4Eg4IPxJkidvDT1KfpOiEdfkZsrHY/KG237p6EoNX9rBcLTblqxLJlwg7eAG82PndifnD
/N88CzfixjHG1UU6vQgbWOZ2FyUt8S44KhsUn76LYjTxUKTWef08tYBU6YitbhTyHfSBJG31UxqJ
FRdIqqMcgUEBCeLEmsJX2gN+xntOzCyqvFGJTv+6fpDpRIkXNh4sZJylWf0Dre7H32a8GoK2n9oZ
4v5nTVTWFPz0pRsxywDUrc0X3SqwYiTY6BohjkHw0MB4mV99LZ7Ut12S5yW5UMnGelc2UoXFHwFK
Ls7FI7xNb4wXgAuVmIzpmZ/wb/h5RFwgiH9I57lptO9aGLSJPtUywAIoLGgi3GmWhFyvzWZU3Gl4
ikg6zodXpLF0PhT+ctbCVf+a3s0whG23IDVM3eYlz0LJHybJf94HoT+0jbOqODucX7n82tzwzeC5
bENinp3Ku7V2/WXS717Lg54m96dEWOdiD8P3bUpfOrqQxNqiJQtVkbSBXwlv7FSIX5uTRgzWmrT5
D6KpnjW1ALv+GNBIqPlxHfs9S12HuaVijPnt8Q/tenMjFUuhJR/SIPIdWjCdIR8lf3UIadx4WD0O
1l+uvhNw1fWOyDJ8OFnqyjR0hqvUaA7XTOyFhNVQ0urAMIOE+tJmD75LuHGGX0BZDJpENOt+31vG
m2IgB+QACPpkIw288OcNDC9Oij4hys0qOaYWOI4gSbxpjnU0jXqtbQPQPchVamCZAoNvPRavfpBs
e/K4ER6rgOTGwxyV3tCecWmq3BD6N8yCh29EEusF//Z6CItGeNdy6lLOFMnXWIA0K2yEt1tv2giR
634uBds+Ba/stH7xfw98qZIbDhJ1x48E1PRJbEvVujlsWNZwXwpdXoyq1tFyOQ9HqlyyvEbXFzIU
S3cW2XVcBNoXML/tf4Jm0stBrPiy72DrBFuK4IhmPNCOa9xjoZ9KxJgFh6eWkhVuQMvILm1CVqj/
HWhcLVnAmQz5aSdzlK8jBzNkzTY3czbPf1DBZlPKAxFQSS3xqGTqiPxPiKa+h2RX/WVpDvK8Fd1c
VUhJF1Bpg3QBTNSH2Mwyz0nyN+6K1MZ9Az75fJWDAAVOqmJh5QqQ60cFMIVtxEB/fKELeboLrFro
RMT5QWG5FZY3UBFOmoszXw4GFXN8jTcX27pBSlt2WkMapDKQ2ZmH7ViO9PsC2p0gUaQVBcq5g1Wj
Qew8RI+SeetZnp4nUrgakPGBfT64OqjfUGsJnDukQu1Xk2s05n1BuI4WONlc1/f9Xzl4EoMifIhV
4fSSqKbHtfn2ve7nw3SEgtQUq7B7pdfmysmca+hi63WVG5vnPC/f0MqVglejDprHKOPWvzwFGeOs
1ug+t622uzVFH7OvQOYRAPMbQFiD2tHEnHGT5jo1wKfqh7R4/nzF8jVugRLf5GDG87UIoXK8eJf1
GT9J88c6WpRcDWwR1BE9XPlzAH/9EnVqbMuOoO/9UnEhu86ZPZwEPbtkgTvNUVf82pnmYv/F6Mr5
3DAX8xvHFIioRRnBj2U19gee9FeLYXXonh8HRLH2fXFE7mrAisZa5qMmQ22lcL49mcAYm+hzaBZA
nQj3Imr40tfb/iewBXSoAkQ0JfMDZMG/dUOiEaJ3bg85wsZE+NHM/OEzsgwVXGP37qr7h40uJOHQ
JrJQ9PWvgKdP0KE9Bu2dzGcNursCL7QLB7Hw6pbyOtfDa+k63TevEgByETNK6e8cDnjSvzhAuppn
HQhi9ZODWMpsbFB1WzXY3elcEq2R932u90T7UJnQjTVCdexXGX7IBXnt9fgMa6uA0nrdjHe+CbHd
OsOGcc6SyKSrgIva5N08HsWeiaXDjPkaMm3/89ysgH390EZEYSTXyMdNiYkW+zY3BC39kTIxX0AY
3Tf/BWg9AZ7Bbqatxtc7HtmdJlBe3Od8vmJIL28XdSb8/MgBk/veERQ9KiWTmD8vIEao6Fyaf/A1
GzX2cG1sykHnUZnVtUfekN+3jIWhmQClZRvaQqKO7spbB778RHz/uYv9wd6ImPs5UzceLGM6NmEq
0dtA55n1YWOKFcADbWcvpTTlZsmTuZ9p6TEY8NNk+xlNSUFypIRPsJz99gFgjiJoYZygymsIabXo
u22+WPbwL4eoWQ9iUPZMWCHG3LfmX1TBbdzElhACZ7wlEJTw+zu0SeT3hkUiRoWCU9y8sPAN6AjL
Tv8G3l1hdapjapjPxasQNrGmJuRnFx3+lQzwgR3f9kJWO0k0z7aB3hUu5uum3xqrONHBqVHkYZL+
zBFRENDxvrQEDx0AYbNx9HHXnh9XJD2j1/aAaAklsbaGMr59SiqkjTO7PXyPSkiYjk8mr+m0/d0G
gz7P6bIW2iF8TNPxB+ohCBr9Bp4wgkfyvrd2eH9EOlxsw2d/l3fV2xXKfufmYzhhOt/8Vv7B5mGH
m+bRoYEvClf34DcPIADk3uBIUShpaTc4Xf3ujcbQg2/6qrQ6rXXbc4BfuFFKBujT4IcrjPRRhsWC
CcWRpYcL7G0vMzf2cFJ+QpjUKb4olhUYPes+wkl3HuhSTWyCFnsaSV4OJY4I6hrV3J2TpbGPZ0k2
+9Imy/UKgtYmENL2/Ef0gGcigElAaL8ELb/Rwql5tvUl05qtw1QNu+SpmIp1Aqif9Gb+uN4P/Jp5
Zy542QGxWdzrKl5D36fovryfO6K7AUDiLryVVBlKxWgFgoM9Za+GRO/PYfAIrfGACk0dAqfqvDFQ
D+wVlIsON9mjnsB1ZJtX5mrYlUwLSaOuZfm/wBDImzvPc1iWiAhwj966Mvgwg/9M0ABnUAuvGQV6
cbn6YAvfb8qskIbYlM637dTAPsQJd2bLqwqmnrgCHwUwQI2RevUdbtuY9zDiEs+R4iQGC/e2mxkS
iu4oxIXs9jx2nt83kSTPLka/AK1Duz+R17P3SdhZrpUDTxskwJcEmESBCy2gHH9x2UM0OVHgsup1
MjInc7XG6EdJmhjqP+/hC/djJZ8S4UC7lhmvXA+38AntIkgkJAf4UaAm8md4Wd9eEZGBaCPkSP4G
uxE+ZQmQ19wWJJnAyaGeDrf4YIhShhn1tMj4b5UVqvnALBG2TxpasxTU+SVeR+dJzw7yDV30kRZ5
hpQwdyNZpxZTj0mC0PgsyEJ21TbF0d20u83Zihw/xHkEF3fOD9w3pzEiT7tTtRMBH9pknlEegv2u
Za+6DSLCV/Ku8v7i+wP+yzrTAtXJvTOSf0gmGxQT3fbTea6o34sV0yXhbKbN8Qn0FjCpEbGNwZXQ
kQMYcKCxH/vezqGS8w23EYueKP9oPO+dN1PS8JgTXhWBD4BBc6KFJCVIsxQI5ds6GpeZtKO9MHjq
dYMJLJ6pOC0/0cR3oruhpsI+HJLGUoU2te7eS86FwbsS+i/qPI+pGZwcYg7rZB7udhAFuqi1O3RB
Ibmjs3p8mwVdgrxcJdXKhAr843ak+eattpHQoYmaK+/oOWoDW5d7YGwxt6O6ScvlbR2zM+3YXk43
7KzqdiCxWlmaOWowI/VKG75jj4qLNrM33rpw4sh34XloTDnedR5xUPXLsYqv8HwfMonlth8eG+I/
v6EbKLn6fpe0/ICkxSxdUZyap4QQmYT54n+WfVn8qzaWUDS9WxltphMwoXJwx+zHwZy0A7FqjQpd
J/LY6zH4xlhCdcnOGbYkqe0Kaq5ibHRdokas9ed2XNznZHxb3hvBcBqI8tvxLXkrk7f/D3JY8D1G
64WuRCJtRpvC/r1oH3w2M5jlYDetYl7BjUGCw1T34jiAWMQ5W/qZAu/hAPg0Yj51497MoBi1d+dd
8fxHbQ8ZOTeC6FVllcTgVB73Gpr5YkOtCP9/5saWJbxtTlx78yjmtTQ1sl96Cdl8cqkEaKaZklF+
6PMS1YqlWyEfdNl3JQ+RzMjhQyteo15sVZKiIGJvn/OfER8TkC3qtR/ziksN6fMMJ4mGtINzNGEe
Jg9qP/hm01Vh1QCkia2gNSLqkpgGEYxtEHpvL5hKfWpx042STyvpoYKyY5dI0RtQD9nIdWTEWH2H
320cLAheXINg7X6OVCtwW1bw2TenzglNZQRiQvK0pLvqbpdilT/6vmtjhTl+3P/QiwYwJFczrFWz
tQcCKkCHZyNWP0lESWHNydUL3lGkOavp8vGsxrCwvO0UM+bgg//K3mxkAuFyy1SxVWFTZcwMdbKy
ac/8Al7F7XyPgnCzR8anP3nq+hby5RRJUUyrOuyGAAEJDmU3coWoYres7Jfo2QopwwLdo4gaHzd+
dHc7HtkD66sgCvofG3L0O2TinoegzJQrErgM1GDypq1a9PUaeB2O5W307scYXI0Yf4/55Dh3SsTg
5nEz2MqXV2BY69NWdXJ0MwloRlZmjyCtEw00BtxgGhf63IyntRSHaIWWZYXU5XceZzd3NdmWuDds
v76Zenqz6GkdvCJTo2SssqZ+tPUMuPsz6dgKzQL2J0QzDM4oRQYHZE1ygK/2R6PNQRtlU29su1LS
OH3sYwgEYVx4pWB1SnqtywL1x4HrreQo88LMeT5vWeQ45gF4QvogWeeC/S+0Sa254+vRxkUe7Cdt
/GPe3886PY8W6v40oNeVCz7es6eYoElbDtjkNnzUwfCt2/U8BL4ZOU8lNH9oMpbjONr8+wNMWbxb
JGCXg+LJzCMdBtkeW/4WyGWKTATFnN1Pll+wEiSv97o196Ha2ZJRAKakC1BWv/0fTZUifMz6GMRs
XJOR003WVuTiAPIjR+U/sBS59qNj15HVIKGQINgMdCBkpWdVeBc3zIsf4tjPVuWcaFWp2l/2yY6G
rp/J7p5W3h6C1+tTYh8AvHZDPhgU8vues/AAqhgK/al/5bG0Z5pQbmMOSiT/xhVD1ix0wbOFmJqO
1VwLTJHsqrfD/EXtnv446374UfRxfjN2BAoA2SCt49yJG2guruU3W26cIsOdw/82ekQQqdE9XhUu
bOLULrv7QiWK+r5C9EpmH9siHNF/Vtkuwkq8Ukc0CMzSrdPVe2nG+JA7LhfV4iP77vz67yLmcUQc
fTdVq5zvqTtYq2b0ALx9fBiA0Rhw73uC3O6QGZ4bpYfmyB6EJ5qOKx1ytdG3ODXM3S3KdPLnn3kU
rAyeFiNzHkS91U0XxWeKogZFjieyh+F5Dd1Uza0E61LCb0yBuQuy6qkrRZYn/wvkXbNfXDWLcS/0
ATHhF7Nq4HQkEG/TtPSG56cWe3qmklNi84UYkxv0muJH21+a3OdRVY+3fwM1LbgtLGxiI27c2XQD
nYBLjvi6QeoN+ujOK1hUEYn0tnw5Mg8mG99B2jEqJ/J8prdaW5OlXm+nc1+cMTsc295LzVAwosWE
QW0iZTJgCebl0bBAdDAg5sZYwxrX1fAIxMH0lvRRspOORFvWToglARdYRwyID27ev4gAzWQGStY7
YpnABm4eDkamMSwH1suBmSpBhMc2bj7c/baeeiHiPzPaeOgR6DnzmjbwFTsV0xpzCbNY6kwETzwk
jcWKiUpE9cr2JMO+MnBOzrKPVeOtSmS0JyzUjn7uDE0MdTPsJ3bMRZsMaZXTkgLZHkcuPs1rr4nv
/jWmKQGQT+xxmb2x71AvT2HR66WQtgStd/oPv8qxp4MbT+ErBHWdBpViDqFZNWZE2NbkwHWk6i7Y
QiC2jeSvXT6hYKf0iPtvH43BLYy3zeeds9WPrAO8rQd1+G/3V+vMWctVS75Ww0xmUx7HdIQK+SoR
Qm4Nfu361iJIhJjRf/STF/m5hj5+abcs/6N/w+u7X33jzX/Ve6yP6heS1VR5cd3sLj0OvrUGLbCR
rWw23mqGzS+vs6wUavhmeMNDfERONaMm2bx5sk5COurbdlUa/Y648SaMXWG9S49Ja5adFWBgyQ9M
W187oMjbQ0s66YdmhfgOILkd7u/IbUVxDFLDIbqhYlgH3RGTpvQ+GWMcMGkUzCBuYxGd5MjGbK8y
1tb6NkgbFQGO8k5w+29pfhAtZO8d327t1+DSOA3a9Je7H4nRVZwOAvbMYX19EqKnKDzeJRfuriN3
CSljevvU7uPHKtjdrSaP51VXl62wwZuRu6IV3j5dhX+IXL06Oc1VZqOLuFs1V6ohljCQfbhn/GCa
2MkzCvspwMzGlCTKHu4yAB0GCgR248I8OAAStbpbJkkNM4BLokS86yh2koxRBLwW+rxipPbmZUL/
6+7U21/tm2mhVFZqtg+Y5oxRRVCI1UIvmYKX0/1VtKfmcjGIo4+wLJjLm8Bcx7MvGTEdR6NO5iz3
xedYnDBp9SRzTlKO60LN6crYrCUQjT7B32UIqOS0f1UG22cHjyM0aawDk/Vc7LukLnml1n44Q9Lu
S7G6lJkHRPvV1AYdfLOvEwA1U4JFR6dRA9g76k0cR9Jxnsl0OGyrBQbgautNmpba4w94898pEyBR
eE9tHo5+OnZKUMNFlDQWJ7ZjLGHD+b59dGoK9ndPuZohyFj1D3EaRiSGjMcPyNWW47ZAEEfOHIet
l0+cOtJlYBYi/d6AFSmG1+cWP+gw13gFH6vWMN2AXctU6rO1uKNNQCjLLbkIDnwJZ7QpsnU4Y82F
syorKeBfp7r+c444rvfToSEQ/mBko5QYo9lLep1/dJX7yNnACdwt9bTzbk6z3m02Zh12DWnmSc+3
s5c9Xb/JUhJl5X39MFzBEirsYZ+LEpNnSf/0UfESkeG/dJEE/1SJoE8lyatGI8x/9ccrkl89tgos
hLidvJsQkiSQoSbABK/H/7CBYU9ck3AYZd4QWWfmQQxYhH7wdGIAQKAUTd6jZuIJ1qNSsajJlmLe
wRCYk85W5e8Sk0D2tD6eSeXyPXM/PCLPS023yc29TNPxaDcLIKBwHIUkhL5Y7nulgvGO9tk5rXSU
A0uEUDujxetS6OUCgMBuiULe+6AIF83nLaUEMEBnSyKGslvEfJ9AGta215e7L+aEkgNR2B4x89HY
aq/KKghrTkLw06l4mMKTSvn3Fu5NcQ6/La8+Z2vjJoPokSZUdNhxeJasYM3wL783bOx02kUwnDg0
b67HZdKo3ukE/JDQnw/zCU3RQk66kDVk1XD3ISpc5lhoDHiCIq0zSjvf9lF1Nnr7adzYoo+87wzl
fM2y3FAzFMrG1CXDrb873H7gifJAPN0/tSAi14RkCRPp3HGPcmvXcHrqdjrBJM6UdJ/Z1W+ECmXf
gv2mByivRofB4Kkk2T2uYPKqKAiIhPrRHERXmNCACqePiTTEo6w0KQzD917e2/deyoMFqoCC/yx1
SSdO3fWv8HHThZzSCmWZ3t07uGZv+x9p9fgxtD08uZGfTco34Li0teXTX8ZawWA3Qil7OI8PxTOh
/PFQvkCMu99uN8stHSCIf00rxL5lriRRtpz2m4B7oKnm9Tr6zLbskLQ2uPJZE/Z7WjC5OwK2i5W5
jBNu7RiNQcVXjo6yv0AbftIYeb+mI8sML32L4H74OvjT2LvnGSBaqJUj+NwKJNBvZO5VqRT4Sa74
VpKFE0BksIUKNWa950/LCjTHndr4fU2SUoSswsG8MySrwwNcD+JvJHO43w5e7MaoFd6mH8wyyfpj
zoIfDMNKic0Z+hpkQKidR04xbV29K7J9NEQKbGIa8ZBKx0/NA64asw6zfEIRSQ4owjany0kl1MXK
Php5pT1tN5dexp419k1+FYSBZEWIfx7IZqkNm43WMlcZ+yroEzl2fpTVtZpFm7COUo+B/G3B6zjD
sssOW7enHRWBCaFX02gSucKkrqFy4RP9kqCV9jipB1SvwDJbC3Xxyv/080KFd9LWhGLScLJtC6iN
TgXOdAXPqJj6jqegC5CjRCkLOy/x/Kqv1/KlwyFwV+AC09HRSM3397JbDI8nKWeqUJfs8PkHCzIG
5/orG4fWCEhcg06p13Z4wTody9hyn/1LsVeFdrxid/Hx0uZTYPE/bE25xGFYr1tSgJVdJt9ZIoOM
fPAPG74ADX//0pg54mq06aPtLN7mJHXiRY1KN9WV5AZHvi181HCeERJjXvkpAPacDa/Gw1bSWCNO
fQFX9isQcnt7oSCHyrDobg2r+wlqvcjZEYX4u0U7aBOkYlOnnOZOB6oH19HR/SEO5n4hHOBmHcj4
2pF6C/iuV4V9H3wd90sIDy7WjlyqWcIMm5wfl+n2ZtOt47BxRwvT6H72uYIVZIFnSQXV6CSKbw6o
lLtBA7hmUXjLzU9j6b/xDTOGeTxx2wwO7TgAhRLsv9gOPabFS5sLRqylbfiByKZLiEOwqkaeTceZ
82xAWpPMSHnVi4G9UFPEtMKzbEBqtzyy5N35jMgkK6DwOUrGj5tyOtcUF53vhKRGdgaMm6u5TDrb
jWT3VBe9JtcZr3nMF8FeE76rldLGItAGMr3CyO4cS+IXyNtR4FE7GKQtnXjCjL8MeU0nU0ePLwMy
QfJptwmaUKELeBdDAaqQWVSJQgLl2XxwaY8HfWJaaMvfT0i/Pp0kzbkED7Dd1auvJz6EmhFWq6NA
GyIkBUa9l6xtM3XzdgKiO68RTvHcA/i7ytlANMwPbnkArzrvCrAW3MNzQ50D3iVa05gaMGg6nZS1
bTpEcqXW5tL96ClwT5VQyMeaaUpTwplU7Z08TS6Qp84iJWLRiIA0ewwhCUYHfgniImWBuNumpOyV
6xny21EEstYaRuwDHXqYk/ZTxTDsFL0DRycTVO4WHbN24FKXCVo+PP7pYt5z1Bv8o6bbqj+kkRQl
Y75Y5Lp37oRrOS2X8hq4H7p7qKIQAkhGQRM5zab745PCPGbQdF9FdzqYI7V7eq5JZkcVhVO+1DJB
8UOJOabqK2L7KFkW7YiCsTJWv7nuwioyk2heWHiMutsd7JQunf8iryLElUiWT289htUrQw6obTBh
ZPlwPIIG2yVXU4K1Uw9q+zEK9lk2hT7s6GNc9Yxze5F1T/FskLx6LJvjN1+kq0TFVWuZTxrqfV4g
wkYwkVxIkCkfhBT1beezVB3wkJ50jLMsWE7g9RZ7bpfkU9W0i2TzWdXW301Yth24qXjcgdtwxyKh
pL3dqPLXmHE+QyVEkWWxzeIOe0KeXsclV2un7EL8WoGkPgetsS6mSs2BFPE6A8t9tu/0yeFlv0sn
92EBoFmTf7G0mHqkRbDc+5T9eVImN5Mkk8S1C/XWEyfgJY0pT0ExfOfs42Pl7JYUvRXUPRl589WW
sisXcoStvYxQQeycUVJ1sQ+VeBynT3R9qocLBLvCc7TGd9WGlfJq1Dg9tR94PTkZo7vTFqVKoM80
o05wHLnMAh4q1SRHLb59T6xjA/bz7ghFMbBl7oOwMHcXhKcnVg7n948mhRnHsaZXuqsJjsg1xMsr
ty8fc7buxvU2K3LDJhVcyIrQzC5zEeLKWfwB2os4a1VmVgUYF2mIZwyMfLSc7cjA+UJg6A2lZYCI
bVTlMpEqkH/QGY4V2nAV8pkO3oIljMUPFS/j84d38OvdDiJP9Z8JCnFJphD/ptMZaF8BIsQpBfBY
1/E1/voZ7mX7n6fdaqHaWA7d2vvuVvY6RQnl2hMCQXS/WRRPItOHIRsbkFHAI6U1iRl1PYT0HLKs
ZUn0RCjP1YB+39B3ySPkYOwJqfKm949lWT2x/xzSy3T/ft7bIE1qREeh5lX9HFU8GPkwCCqsoRBk
+6154S6nJA5VANhabG67AXQG0whRquge7/KZh2ZFn+m/3xpQl9K8yAme5c/0ufslYGmPC9me5CNh
aeTHBFR9AVtaka+wt7jlw1+HLQ0efUJ3CXiQW5N+Oj3AeKJIIQMWuviMDrQpmpHgKQfRGhkdDexo
57KVtm2DdO/xbMzKHCTV+CzSfw+THNpisDgpLEEQPfDNY8r7EN18ToG8BrimJ8z9EGV3N/q3/0sB
pphvq1QtfbX9mCy9bmh4so2wpyrykw+urhb7H3ubreQsIcAjcspAmCcIP15ba6vylZZyY0UR/kEF
xWhq9jZkH02yeom/ONf6oDQZXth0BXNmhWC59/3MLjP+rHQvT2M3Is+OeR9IKhcCptDa8GIJ4T3q
90YFO7VT4reeVA//cb7QOONnpg4QrlmjqR6PIMCWeorK8M7XB7/RTHascvQCzJSfu3XBeK26LqWI
HglnQbj5SPWqGKdqdICypkzpx8ajIhunIHbJPcplqcdt2pjuoyC5PUXJL9Ow6JH2tKX4uUPpAne9
KEK5y61r32tVjshiMyOVfvMflZfZVpr+JwRK3tBIplZN12nPwwNMkljbyVZepVei/AjMSx59eWnE
NqHMn3CZDcolb06QSZ+kZjjvAr/qrxKGTjvuIFndyMjr45HqIDCcNdzrzfpzBKpPIt9ATyYRKKnJ
OreYQlduINyYHePdUP3tC6Ae/v2UHG6Gidz2/ljMi3NJgprtkKi2pMyZs7ImXFBMTs/ZkZ7XDSnf
AayRMbxqYdQUVVE794aTDEz7m9xYDsdnSEydZkxpVOVYNCLfviitInBEwYC/t+05O7tbo+vSHIUB
4iFHlQxgSkXEWXzTKtqPrmP9G4V3oDK3D7X+Z8A1LAlU6JEaKZJqmar0XrrsRSYTOQZ3GgBWYI+Q
LwZf608CDutcQ6g7fODzuIbiQyzpG/dAPgEbG/BGUhfK1HDN1oWzTn+ylB5YkUinqdKpsGHNYR5R
BkcmCQO8ZPol0lPB0wVm3heMlqqtNYms97HuAd2uMEiD+5Mwn4VIgWkTyySnXO6WXmESi9FGfOl6
fwA5k9uBZnDt5ltR2+DaC9V9+Z8TMDGo78BkQkR1gwQaLBAlfzLqmHpx3JrJbqmUh+8v2UZmZjWM
/nYphfedd/oD5UxMaeyP7BSWJ10NEORlUsPhTax+DT3CWUkWrKrH3ucYTRBYfHEOpioKvsZFM9UN
3yi0z8DjwFvb7Lso8RVclPd7GmpiG9dQKwphP+E9GoUZPO4mny8UzxCTt2vNGUgFWx+BGm6o73t2
erkoAbFszT0ELdhFiVOszoCWK0uF2dz7tAGXia7dswMRuaM1JXOE6hCfYQnHcT9DhKRX+0fLnGrJ
tTCCHhiRqKJiY89k33aVFTeBGlaQcfc7VmSYE/Eo3EvkdxBKWoIs5eFOqcFP4rEDDLNRsK0DZZ2X
4BBON4BgLmAgaEhxf0nO0P1QpEEDq9S+QpvB18nqZQ8mslkVULVLEGvmMs6ADYv21qP8Gw2ltO5I
Yoi4Gm1MW4wUlcS7ldmjE5dSutJVw7pcNkNvrtzreyg3UZ/r3RFk8wNyRG5VQWiZeenVhach/PtC
QZFaRYXTxgo/NmRJQbJVkYNCyVXce2dhJRvvgZSkBxjM5OuuaqJd9WHFRuzf2MAoKPJ6Xi66Fdlm
glLBmTUq2FwlzhSmCx++/k8GYThC70eY/BcI8fvqRJsz211P6zzQQHsGfqh6IiGLuCgWh2HiHE7K
Y3llpB0ucgQ0WugYgbTElLdS2oAFM6ubffdKAERjcxHufv7ySLsyl28cloTQNcz/gMsZqWtVqIdK
AaQCCiQQ6xZYy+1X26Ta2rE3yWpdTebJnRuGU81eH1ipzsz04+L4vnb7LyldCH8fAU98GbN66y2n
uBSYb07aPVvtt6aW6HYM1GgYd5haI1qtLtOPnlZK2UraBAnEwRpVz+jCbLaKsqB7K7CLvPJuctTd
9OTKkHApvr9+FL8VskBS5yLJTYxYq21Zqzazkb0wH0pEadjpMc7lC5vJVFcFOFLS3osR/UUa/ycV
C7VG7R7hd6wB1X7cC+ELnUpFh4MyBu2l2B6IHuU4iW7nzuQ9lwatqbSi0KgAu3KkP4WlxaWsItuH
S6+uPkMmkWtL7vNWhY2BWBR9mv/vpOM+BFQ8KMsNIa8SElAj3QlWJ9ejNkhoQN6nF9cXHauYTzK5
uNXVIk8joZjw4E/DZqpwUN7tTCiNFQGpR/1Lx9zXixTxkMX6FSP2KC+qOcuQvmiglbXkW6lUkRwj
OcyJV7cF19nDT3tPf8UVmGl8BBpWnYudpYmsB7EJCSTtriaraqCXj4fIAprYaREoAD9qVRyytAQx
bFp966VN6RG/uPv+3Phpe5APJxfdkM5+D8zNOoU2C/GWAX9J14qMPhtzR9+NKxfH2fY+LWRyZpji
Tde2xYMCxxynJRqcGe3Cvn5gQ8DTaC81lX2fuT1xxFcLAC8Ca38jCV8zeCauG3zFIHWFCLNLHYyH
84F+m5ox0Nrb7T3gUPz02n3zutWr0QqpnNPMib+6x7aBljV7REAEw/rvy9/Skl0T87O3FpLry6Gu
ZY3/TksooFgeOy8mGk5xcXthu0zn6+V4SlgW23Re2NmFJrSgt9luPjj5ANMIGVnjzK54OAFSQIkv
hBGzOt3TSn6HWPWaKxpCYi90uzx53XcojqF3dVg86AtXnr679fhpvDqnHmdz8lQJIsIK1+sk9qCO
OSbxjBOVQFdojp6UsCRKWjzhq4exHO5iOIL8Xkdc5Zv6+Iq6lzt5e0Q7JJ80/6X6yDTENCpmu1fJ
7sedYaZwhGnRp4gwmDYey4A9wEUhDnRuMk98mGEtB6R4KtmO8fOx96LIJtICwM4Y0jRJ3dXw4Xm3
jTURGZTCQAn1oG+iLbDzgAjExM7lz2ppDD83ADUytvFEc1fpAGuzfrhgfzTPiw946twuQRlh7ASR
148X+FImMdxYbQVpwJCBIm0DSwBEE3atN9VazZ5ecBan7U+z+JlHT4DzKVwTLpLT1b/cjkSChRsU
Kt53+SWhTpjC/WdPHNJXoACApr9Y+JUgOJnrG81WgFPbaWkdeQLGq+pLDM9eAi3iwA/K+PpNj2bp
RPAEb0pk3Ytqd64bQBBsQXWn5avC3EW5zSmdw8ThhxTwtm4g8L0gnd3Q42tF1zzbcFKhQ1qOxqlY
yP0UyRRrZs2wfoXyYT1ez0MFrWnscoql59XPRXnqxCJ9EBKUODIDAX89FTvWjAfPfiMRcK/6jA6K
DgiAbvTsQO7f5xf0SI4v4tAvQTD2KMO9Gb3Y1Rh2oSnpmTJ23LMfJl9kGP+9Y2LLahkjFURGHzdE
0AGqU+npYLv7P6HAmHgH6+QWMzVi7dqjYL4FE6PyHZQRF8aqIeodUaqawTVtI9wFoynRkuL7gyCk
0DcLAIDieToxox9mWqP9pm6VHetU+zDOX8Tkj6D/GaKFun6uDswz0G5/RRfp5RZACEb4EFfR3dbh
39mq9R52T9BSOHJXBoL7yEKVl3xoWivwYXx1ychmbecNGWlZrgD0Qs/7STYfZUna2oQEK00GPw7T
OatVVqUWSsgdUF0Z4CAYn5MZXW7Ug4uXisyxG+UZndRnEsXoWcyHg5DR0HCNunzWsHChfTBbRu5g
TmWOiePnbjKvMhOLh9TCT2Rgbnu/SfOv56S7UFKBJc8Oz96M6JtG+jIMuAE7sDZJavHWZgG0QHwN
K5rr9G0Utr7+zOUfO4w7inZplJL52npmbS27J41u301p0Dz5mxD8HNrfR6GpFxDSczr8ENzuomk6
/JtTVwH/EeS7bEjTjJzCQpaOaPAG7eVIe+Wt0li2k5D7W/u6J3X9BGSSN5JlQUp5JY9N9Ux1IBwC
kMM/dwxfnoQ7eAcuqujAwTzKN2wP2Ew7MA82KCOD66f70HUEHbuODO6tmdKwV0C3ftXONnLqBasR
dHvyDNO/LxyZjgtzOUW2Zkbh4Sv9Deq2J4lEt54Oifc0imy7LKAFOdBZvi5qkF/aQwrf1TQvpcQN
itA+PgqKOx1fs/ji6gARy1SOnlDjTP0rhRP9bByBHp5lzbFeNXSjHdlcB6u/ai4eS+utaTzXDiLG
yBNHddyJcinyW8Eq5+JUEM08+PPf78iQdk8wxsAzI/9iDfzThfyqwWycho7UBICsrIdkI8TrEfjJ
rqrUiDXqkf8r6Dgog5TJl7ifJWnG+xrELY4UlVXbTYWJo5EkZJBkzdNwBN6bZzr3f9Enq78l+aDs
SyeBhlZJLUQ3nOSNNiRYdD+l5MJJwFSQewq77qxk/YVsT+G9+yfMtmec03DTYclkUiSV5eA7a7LF
Z+qdY0qw0ljOrQob9TBj1yb6yzASlG0OA9EA5Td6GwQPElPNcJ9tsB3T+C9kncm9tVTo563wUlZ9
hqBoMUem3i7UFCacQT8Tw0MOs4rZTHjG6KPDiKv7k9oRiBmnegYpRuB/LD96FptgQU+87jF9I0Hz
sjUpv25oGRA/lYk+eFItZELp+r7NV49CH6jA9W3/tIte5tOMTS7AJqowWsfqTYNifwloB+YaVStX
eMMa/WzjiHbXSSXRbIV08pX8eWyl/wpc1l6QV8esKdXc9q42tfCEWWzVP9Spnoy77XkxKWV7Xl55
iaH9KbpBJAL6Nf2fuo5bZ7GwRLre9rwe4Wg3dbUkDXw29wA+F3vnMa1qrtfPkVQBnhAB0X/C66b5
k8XdKVzKXsM1mKEb7YVa25aS14UqbwbLM4GBBKks5vOdeXb86i8l0fgNAtGevn1Z8SC2xQDz5Mz1
H1EBAcbOcUz/TD4NLnrUmAFMuQ7/7Svhc+uCNEN1SaKJs31i6QC0w/dNnQogqdhlMODM5TSLZszb
CgBB2yUgpj6kFVfd+4Ex5/tceWjH0L4mfFz2j7zlLObCg/EWR/PodpTyTh361Dkyeb5I4QxZDqy2
gcJXc1sU6C8Ff+AG26des7TdFNI0MO6dH4jlf8ti+0wWSZgQEg6qhzhfqBMCll8wW5yKpX2QBpny
F/xgeNz0cIKd9cF6OK4/RncW3jxbTAnzp0KkzyFAcJLKYYJZjSnIbCerWFiKBZKxv7c7VXTHjGji
ksYxyYvPV3QAU07LKr2zkjqo7/ylAC3QEKA+VG7Ra5KXYpb8Kh2NDSL9MJacNRRr30zPnl0ytsPj
+gS89O6N1G+ET47ICxlCM42AjINuZ4IJLqPzyDw2geG0xrX0mWXP0f28qGAmRjO6DSEJDjnkAL/s
C6pwkzwNZmvbZMJaNFS+zkl2ePDvYRaEccA4Xiu8PS3kH7T+F/4bxAhIFyPdp1U6tyTDWW6HET5f
v6AazvnP4vMj/sAMawXk0Xg4xuW2FMFYLlqyXl0uOoNXF9BngG3JqaV9vXcaoE7CKtURjJzTP1C0
l3/7TR43zRtomOIXx6GUwmGf3AOgwKe40JUtx7584K8hJtOLDqaTsRgB/G7yYl1CR4AnoC+4w4yM
DwotCeNvDmh9Ceeq4TtmcNcwM907pQSOg8zsybIScK1lt5nrBPTjJ9y1MTBxqqgVANUEjJwg8ua+
HmZjPi/Yf/XdhUxEatWcj+Doo4E8A6M2KTn00+ts/iNa1p/rR7vuPcVOcdCZSZkAvxdTr8b+Xngp
3wV+jvZ5BS1boGejsDvJ6i77DEL7YrYFqJLCLAGZ+yaHxX2uV5Hk5XgD1tRpf/0O8LpdWg1LXcIg
qVSCudibxvQlsVhLusqJ17Ta0Bw+QiozSh/BOgTiuD66z8dqmMMKqSuP8hpQakHeEZ4H03+oDsRW
b9fZa+XWgZtTefxwRNr59u3ByVzOs7B5GrBWxF4XAvkJ8EdTkSsFxjZw556udnmmz812a17YGjcc
Jx4DlulhgHF+2gGoVoXx/UhCZwH4tSJQZK1GdRcHrb8i/hxRFD6UooWSLOrzPr8uGgqrYXCyVqNP
3iIgoS5ZhD22LxW1tLipc7PE4cfPf1gt55DliBgFf4V0PNmIo6E9mRd53tcOC4lsiwsLCe5l0Wer
AvwfldIx06nJiewmieAXXzmDSWU5Ska0EAVL06nSNV3Gnk5lb08l+tPPp/ttoukuWPX6v5D2xvw6
mStxQVhIh7WS43P/Jg+ZUnwSmEDZsMJYR7YtGq7UrkHg/3moxPup+8Lc6meCGtCqBUaemZv0rZ4j
JdNNiDcgnXMDApn/0VaC1JL4BUCe0PXOlXhxluzeEi2HVTGFcdTaGQ7Zl4pZI+i24xHm1usbWJqK
SiMVLkc+X5VLHVJDUWIznYpKgL3THh9PzxOfM89NEYBbArMfER1siPv+w+EuNOQBrBi3k73iV+Fc
WGqd/JaCm/zV0MCgQIGWzEWHUH0FuPqxp7h6LwIia6yzNJvox6T74gaWJg6hbi1WRRw1CjXO0n4P
QsKUnlu2VwxSOjvSdzmaVJhd3DesbLwoxk1oOLFzKHkcMliOC9k92NRz0exixDi7Dx9ic/JHfThj
c03ZAMWm/eunC0ril4w7OEBhyN5s9NFpg7hOU9gSt1Iu7Iaizri9QsjgKQqsiQRZy4A2HTofuW87
L0a6uyZKrQpCP1A7OlIxAnOScymWSkoiPGaKc742z+Irot5onpTObqkQ01KN5mFne/6SpDh2SooG
GLN0Ah2YdVOSXh3CE+4Ndz1au0R12gLe4DBShi4qeYYYCsewOx6NnwEc4njOgFVgGLN9/D1AEPQI
HCn0og8ks8wj3dvQoaPbRAFvY6xsLHw3ZFF1pCYYi7y2yjm+414TsBU8AaQaMROcM5eUIN5p/j7f
uMvj9e1zKKNsYTce675bo7fJ8CSx2VHG5GwWWe92KmYUL3jsRTAC6CRfXvbbkocmoeF17zxuOzt3
KlZpHMg6oQNgE/w9zklO/JnQSWxiEr87fTXodKfUvpeQpLZ5aYWoX3OOs/llmM+w8GG06Nzlm0yV
dH2skJgbbMQ/62H0YUPU65rBkGXzW7bRT4jBy0mmfICyUyxNZgmI/Sk5QUX68jygbiGFRR3E8VX6
veKQfTYsA1t1mhzWH6SBFi8oPODTO4b6ziF2rN0IukNg9tcobivxcEMOMFXRq+PnKxEgawwQvkid
M0DYuLf1hJk2yGE7GwebNZ0fBYAC7XplPAy/KilovyepHeFDvFdhQc/ZmvRKeevsHFh5N47gwfZw
+2Xzy2Z0LnqFWlpejxCNdXSpxPHOHbn9Zqlw++XDiO5IgImv3dgc6Qhxm5kvAuEGfQMCY+ii1GTY
RmcDqqhBPiTV+ivZZe/gMDmn+2KqHARUS/zBe+OE2iw1h71G2Exd6jviS2GLA13o6+K3YF+ygl5u
Bx/+QvN+aSCGsoAz9BfNG0WlizE4HrYrtyuOURhc3kMegZZH4cHPOpCXrIlbbwHLri2ZkQfdjQE4
jfppW7GD01jviqUIEgbA4HE8rCG40jwXNQrU2f3jQf+oV6I14I5V2dIJ3+fKJVKTDHG5zPSIpFJN
eLj4Noz1kqoS48VJxEAMpjjb53c64lzH+4cLGeNG5z0ca4toiwjPTzgL3DBGcshNDZuAfz8ympa+
21atSMqTe7NCIHbeLgPbV/ws7ORx/Q3ggjGFf6Kxaao+s6AgF8oBpvmJ6+BHIrX6bCzsq8obQ+mB
mB+T8901c4aJ84S40AYf6W+ZXEi613nhKt8m4ukZw7NtgKD95tEZpRyZzP8/ii4qg7U+n9ahuzt8
1HU4MM2/lij6EhNkxewSyEyKkV31bCyFEw8vMF+RkSwj1LXRHI/mC6B1DDpzoo/2W6+l+A5e1yXq
EvPwFPGsczGJo8a7VK7esb4+PVDAcv/8qRZx7cT9Du+U0OiBKquHmq47UdGhB7fMKyH4WRkR8QjG
T5AKXiX3F9eYXZfUVNl8dAo5nyYRVD4SS/pbEu2rJNdqVB819GalPQyaz08x8vSE6H1KL94P+alQ
oaa4h8a6eKZ2pV5N44wLCIw8Z7A3O6T4qiizxxo4GNKoFSJ0gRaGt+9xLXEfslNJ1NtzEGhQllYG
2trUyWDwDhvsdgwk2nmjNFqhsSXDisgHEHWfHRi1gpxO8nAPPt/U8/714SBmBYSfeeiBe6WViUZV
aCpvQ1BzAxLsoiu3JC8p0JJT8HSXqg+ARncMMEkwU5zcMgw/C1gfNKR0isxIHrGl9G84HoAyyWmN
F/2f1XXAN+KvO9UAFap2dh2206DWCWcR78Ttb9c9Z9yGC5tvdJIPadeHH5R9K9oR8PV7zQwW1aZc
KraL+oBTJLDkinqDJGYJLITlmgaB1lyccGdVcdMXQxYy/onaMGG2nIygthlrvMz1Y/x84qYewYKW
8G/cgrMrGDrkKJrQ/cfybbddm6kshZEruFPt9Perx6HbIgsCtvjOp0T54uiaROzKRQ+8EuJFayJM
IV6r69grZsNhIpBnGbKmthM00d4Kazs6p3SWVOPl/cLo0KfS6goK4zNaoZL+aVDQJoJqI2ZYowPY
Yaltixmq6S5Sg1ZeglmlpANBRlx2JJsLYRoUdTGOKwzM5udzYwBL8Q1H5L4G6SsAqANtoH6kh7mF
Bmu3scD2aRFD1pDAFyTpl4Ymi73i6jkgtOIzLzntXtjOV9tJ56BmX3V1PVelBaT0K2MtonbRdeJt
6QXTYFflb8+Gib7+z7hrCWw2IB+iYufCsM2f+aA/+LGxGwcwSS+hz28TbKsrizgWB/1hWkh9dF7x
Wur4Q580O6i07RDrldWDU6fZWnGGksRlW9C4iYW3tGoijkFReuuGEp3LiCueVrJVyUKZfWYShZHL
C2v18cTIdnpUmJZcKpDs5GKekk4MsSdrJaFgcKSJJI1ik0GJ41Wkeci5gprEt7nDe0+UpJOQ5/qY
5AN6oMq7rvzcGHTkVFOADVXDTfI5d2+gdH78GhSECSw59OU0+lLDa39Cwb4wywBfT6R0PGpK06MZ
nSTGqyWi+g4qXlr0wUltbaO6jOC4TXTYwNdlqwqZSTRyNZyPa5VbQ3PtNwMkOTXdB+Pu45do4obg
EdmPfVp0NOnZaMMGVKhyJ1kyO/OU9ENDDzoS8RdNaEwUIYEne4uGgYGDT+CHy5Q2ZE1KppLurh9E
djVIlux5YXl3bIy0w/vRrNSLzCbiw+OxQ2u9rrP1xDMMZ/XITJMRrE0PBgCkQt6JLN6oSBO4tc8v
muP/M0Y+8ZwOST3s/9JZzjccuhkrMVbSHbQiIKf7iVhU2WGN+HeW3F0TFKeUUK24F0kA8TcVnNKu
N+XLOxOch51b4dkam6vPjZqoaZ7w4hLyM4xkWwIha/X0X8/iKmSDUNitOwRnB+YulOotDfAAp0Qh
bWK9g5dKerd0tjzjgLAD6D/8MzTlKWxWTlbcKlfl65IjSBQa5nFvbUzk2H4BPq4A56YtTMoK4kfQ
1vDDT3s/JcNvLM/MsaM5HZkyY6FtHL/pV36QLcgNOBNMSkgMEqovqSs1j83FvJT6AhlH8RizTiE9
Xyu8FO9wGbgOkxZPM9ZvCvkkpuLfdfSwuNZGT4emhdbE6bygELCogXHC93xL1PiPMRZo9BFa/7Kj
l6lfnbofLqGZFRp8Ju55xcxdIUlj4ahS+mwn7ga4CuIqJp/L90ZRLd4zc2fSTA5ilQcy3Rva5wPe
x79fq7s7WjWT+bYEnJqGMhAgYDhYlT27XBFGIyQXhzGGOZ9UXVEHxyVGuxzVyx22rrbb+yTZjx0j
6ro3vxdf5TxiAl7U0Ob6KKPOKnHGfVUn3zs26ITfyt84Cqux8TSCkGMHf3TdzXv3U99V/VBzXzv+
M2ZG7ahkvM8ni15G3bGwRNn5CQnYYbuq193rBR7Ej29+q3C01A6EY0af1+dNf+Wc/5n/CWWbuUL/
RKhDG56LGoe3ATc47qNLBmiMQ0okhVTpp3EXS7lAAJ6zktNG5MI5QYm4kdgzdGDWKMI3o0+x0UzH
Y5AfdzXmdfFS/1No2TTNt701TtlXCGNZnddyWsGhfmnkW2ict9N3JQ0axJGEt/Q9uEZ5PwUl8jvS
Dgr/vIrKNiD9drCEAbQwmHzTTCWQo/WtsaWnMaO2ROPj871p6evyqxrjZHsVZXsqxDbvcR2aeqm4
bGw7/jU+MwBFxpSj2rqWQTXLl9v9uLdyDlPTZzAW4Jt4DVrpqZ/RLjtJNbfstzsStmA1Tu+qUFzD
x30LFzT10Y3M7Xx64p4mj6iN4LiHGugsnZkh6uCDdKeJoku2pePRA7YxOg2mF3ONRvYvChX0u/Gw
JwYdpT9g2NW5ZDyHkUUCfOO8AJaayFniHrQvrfZC20AG0idE41GFTngT8xoHuwlEytelIUGYGZTQ
DMzjh/3t3Z8IoRycnAIUepjxyRvVipQKIQchGIdgxExy0Ge4bhlBwo88MwmyCB8TXrwNasGjRx7W
Rm8oSk4ZjsNWDy2oa/Ntq/dLiVaX2fKPV4lWh5SaO0ATUWU7j6h03rJGUj/rEZQGkNr1r5LR5YF2
RUvz8P8kL0ZOp3wgBXH+H95chEobovUJPtcJVLFIwFu0hIPB00YTkhh6yccJ9V3JsL/FvNLonz4v
otZjlg80wYGq0m4tWywrRudgVABWWhG+IV0nQctmlVhTjBwqBMRGgN+r6svQF0onmoahktzUjuXB
BZLuFmnnt95LpS9/nBkflEgJz30LZ+UeOHazKhmTIYZtwDRlpG/P5HnYBZ2efKCX3ckaGLKXpJkt
tOBqCyDCVQhRY9mc+fWvxZhFT7TcTItLMM9knP7j8PMuG7FxrzsUcd5+zZ4HL1dzgnDfrvTGQSL/
WtxlOlG2UxDu4B+lcOVfRMbUrsLctssfClc9fasRwfDKp+NZScy6sp3CgDn50iAS/nL4vJmR+qYM
68HZ73xL8XCwXVVWHjSFpo92CWd9y2zqna7EtXVxd22rLJT+5gEnJMLehPHr5TlAHwXkGnX5xruG
3uURWkgRh9vI1kt0BwSxXCKGMj4gocutFkgVm30RmZIFMMYrWmtPBmIZZLGhuznyJjpR/2ijqOGv
I4yWNya/ijUnwUNWdTAW0gO/UtXyrZr+vIti0zvA/9IeCJOuzsnBqRa8q3yaYEd6rTxeXo5bF+5Y
srhxPiYWCJHDt2dmLGQDdDQ60hyyfMIF3taqxwMw1scCPcEWW4ZhsCd3uED2tE10iSnnBzbm1oJH
/dzZb5NxHbn230T33rkN372Fvr2ZkzFgMyv0DDF3iU6H0VpamTj4b583K1j5ZKSL+b/heSNhGde/
ZT/uKUvZLlc97miUwlkIyacW/pbMrDrUl/Ymvbeb3m4zG5lIy7Uu+O4xU81GfZ8NmFV8S6O5LdKY
2OcdeSdD6RzfOuPl4tzzcumMrGs9eih9ylbDD5xTU1S8tZMgxhGskFmNxIdvP78DYcK5xBV03D3g
KGOvaCc6Wk3RzXxPED/QRCGqJwFY9V5uLdEjloiEigaAGiyVzd8vOnTiB5mJYT9LpxVbEFaJV3AW
nIJr97OfbJBkfGQ84nw2VRLgEhqgtSkmDIF5EA2BQSI7+FUHl9H96ouql0kdx8J5h12962HO/suG
0OIljd+mAMavCLf1Uti7g4hcW3UFy0P9BF+TFktfS6RiCXI9xuJL6zr3yUHEI/yXFXlvCp22Nq40
aDPZqGkrJVKzqJ9KpXdecUqVXN5/RCiPWjEdNNkGZrC94w6wZauh96p67MINncP7lz1f2iaAM9yH
/HPR0t6QR6NHDL5TnByZm86f1VTvKTvyiRNG507IwTiDrgJ6msxRPffLrC/L9yX0GpJwXeT6DdGH
GbZVi8BALLynZbSilLPJRw+OQKktj7UGUUSv78Vceti6i0owweC2EjG+N1bPnYiiLUTfDmygAv8U
wxiPxfMVxR0cJOoxlY5rER/MPvuN5dDEuJV0w/iJx3mRHiGzIJRDpykUBLOqnpYGxpE44galztfs
Z/m7/PpHLLq1Ewa4OcIdTe9fF/N7mlO9/MK4jynvSyuoCm+rFTvTOQDnhfT1fEYExKn7AI4X21zg
3pV6DFs+ThLx1QQxAe1ELSa+socm/0xId7NIMRlywr3L1op1reo1sw/1r+qF9Bm/HxhapDJyhumY
ikUCxbK1LoNcHKwuYMPVkzfouj8VmiwBwmsiVFp3QDctUkH3eWin/R69JT+PcC161IkgthdzSuK/
FrxRYq+F+MeQfhaXe0YNMaiIopwxrndMnQ+0kWLlvO361qwKNtGOrS9bS4REEYNlRBB5sYsHSt+K
/BWOTNtG21/aIQwFi7rGaypF891uMIwk3arRB/nJ9Ai8x9OU8sKJnCscdUnsGnY+HDd7FV/8QutV
YXmB+s/Jt9Db7LVNOaTDk5PYHoU6Nc7oi8ILkWa4mcakJD7EuPl305V5SPlqBhhXmGKwZwkgwMb6
96tjiQPbsrEaoUal/wkTJYtosU+ok/8giQ8hjUPYruH1hkCI5gQzH5coLlhwKKxOoAvXMWh0BMAs
ZsdZsrndeR/fEa3CFhjq9J4MQp7vEGnYFEtou4hwaJpza7exyDXn88zWPQMvSwB2lE0N1zBZO+Tb
3XyDAqRV40LhyhRaxcmWCvpkdqXLRH2KtqC10y7TO4dfetWnwsA80j0lMjx8hnQeA1LKIT81yNKj
uGaZ7yNowAWKJczwPHz3vS2DlqLc9JpSgCPxfWhXpfKqXvoxlB9f/+qDc+ZKPGYx09wy0+b4wS1y
xieQHyD2UmetBpNNFs4XENepRcpLYV+xiITSRvb9s3FVQQPXAHW0meqbeSkXtoPaPT/FOUrN6WIC
9dHqJs7zol2XmhhfwLuCELCxH6ZA7To24rewJxLcsiHKFicXgajN/LrqF1HAm+lButDPIBWLFxY7
KYkCzaBuH9w9A4t4Xcn0zltxPVxmpf4EKXm60+bm+apIAZseMZ73wUaHbEy5pS5ivmFkC4qFNuWD
F4GmC5J9ItYiJ5QUwuhp8/HHe2AzKOPlBNbrMLdO8YR0+PgzW++gr2XfloqB0RYG0SNSA9szcEKX
uDgT8rTzwX04PqAjI6aO+44UbfPMuGLoJOfnqH8mQF+F7qtVCYR9ccDoqw4KXNTPv+LX8bdTJtdC
/5GwbjCBHlW/Txi2vQxmOLtDrsHwP98l39c2JoGbbWb4CWnD0Bm2ZujHVLiMAgu7OubnooUcRKSG
agVOJioGrGBQsuXyCJsYV5StsxrLELQPI8ttU4iUOt5rM75Hl2f0WEcr6yBm0NTC90udqgWB7xqO
UJFVovPFIlq4vAE2lCWwj3NdACf1imskVyBSbyg62qIbcW74yKE62Sr95/Yrm9DeIPzcPQ/nfPB3
cfR5TdjfbeVjyPGHw4mBOPhjaFGf1PWk8OBL2sRqVSLX5LQcHl9pCpTNMEhD8YxqpEmjxhZ5U58Y
utf4AWtNHE8L+rjrx1bS5zA6Oem4pkMXUxHCl6J8TDi94JWZvFtSFW0/ULeKalgEJ1WvYtrSn7ti
hibXoH8f2leWV5pJ97vjAc5XJrmxyJtdyMEayNi7RbBlCwOPTctYP3DB3hsGpgoxJlztA2jsOheW
Yq4FSVID03xmcmW7v2Q7p9EUZI0iIv+UpCKsa0KGDVL35igVNwjnCmyn9WatAhBhqkANRKQSbJKa
tBYf42I9l7oUDdW+dVm4vkM0mpmHMUBeoMLdk5Hro8JhJ/mcDf9/Dg4Pd5+/EOnR7RsRbA/Asyim
V2xg8utEMa/C+igQJw0+ZqWJswQiejWos6uNtGAMztbMOK8+enH98jNJyZ2ndnWUMuQhjX+poYrr
nLdoGvK8AZcRttBKBLKWk9LNktiI5gDUb/TNHs1xfb3szC7P3bSsnrH9AltfbSclc84wgZy2iyaq
B8hec1skyHqYwg2Vr+KzskjL/FT6uHJAcbYcXkwW1r8zpuebbFIziIgnC+5c3EnDNfpcCbTPH3E4
faoA2uAQzkmrP2/nC/iPyAyw1HC2pZn7wDEToX69bWfZA6uIfGqjcpGdsjtteBHYfw1iVTCvT8j5
TKKZnkmgfsNdRFcZ5kYxQH8K9AdEZPkXl6au0rKKwab/7gH3qhTXnKoP6pbI+d7Wbjh8KAa1Ww8H
wC29DTRSn8afcgK6+OlujRpSkF52QWGFfSYszSRMvPdhXQtCfyJ+6l1PcTIQOcYJ4znMQvKbC75N
6UIR4SzSjVvnMC0vqEPPk868rzQT3ni++Sb3d9BQnbXE/Q4nAqqs1XGI3ffK/wmlzt/Ca3QfsV7B
KKfUWtose7LYup5G5CSmXAbBiBddVxHnI8EkfQKY8txSDzFxa2U/ViZGhNp3YIb8JZnhYJMtEihr
bTqSpHpTGJUOi2ypCJInjUDiX9SsBdMNHzQb2CJpJOwaPjvYEtTieA9oQeP9RQ3afEOHa3aRgmsy
WixfXQU3dOqb64EumKzZICgULuRyKzzmIVDUj0oYhh4BGIFXvz+3xn/stRaPcd03Pv+YZKb7XKXB
NNrJV84XF77HcWcsxoqTzOoEW/h0V0viZVQX5VkunWUpq7iBeqw7xVmd7IhXgIN6ljDOeF9gUU71
QZj1L3g52StzwLczvD0LDjP4l2zBty3mkr71amOuMu0Dl0qaOr3HZDBfzawmJMXvQ1rzjwbqJGEC
YltRtZWuMI5M18PwUgaFFEVrELONacklNn+Jnjkluw7wR8Vc9vYSOFMoqa/eWR8rFUOn77jHGE27
LZLUo9N0nuRn60YRwe8yh94EAjvw8n/hM5EuKOBBiIfui2/EwBJ/x+p1JOfoXcLpJHGluLVloIkH
t7trs6Q+NwfVdUteVjNp7aAb1viYaF9+hrmE11ZGdlMqYVYWB687dyQvmGhNtXYwM34/BLt3nuaX
agNdrXlruT+ADGK3TSoq4+3T1zJCS4IQU3q/EpijJ39uNv4X1Ruv4/RK4EdpaEFphEeKrZ3rGN5v
xI3jZUp/vDPGD44HtTq69d5SvL0k6hH42q6tsfCjJinyh7AOLSHaPHWF321NyTn4skz2EiXtquLw
gYfStE3/5DqK+W3DTyEPcdhvOFAbIMPTO0DNF+ZzHAxDiOVKH7v/RNfidD+PxERXYTNN59TWxP/k
HrFZC98iET2zxKAfc4DPA8irdqubni8Qu5NhcPW4tlthWKZemstnhtix0sfyeXjj8YSkGRSHYwBL
l4WSd/bIJxHz9ddlXPGdFCyjyv/bXyHw4YDGrGLbM4Jz9WfObt/4ZYhE9hS4/5vmsGshRiQJiEUu
m1SOgvvT01GROy8MHj9CdxhrYJ2Oa8RNziYKPmP463optJv6QVIwQfeMi2YWp168X2/vLbKV0/rK
SNN2jCPNTsS/RNjOdqYyR9R1z+dZUnVZ8pEDJI+1gtiyF+PgTXyr4qGJ7W/M3IEalkkM7h2TpqxW
oaeD91MMaOM9yQSDA0BZ1K0wppYsJXMMpiIddS1UUhCaGny1I1GaaEvsGP41eAr5RDpXddr7eq+X
mQh4Ptuyin4uXTNWN3x3KUQyMfrzEtV8FdS+VLPsXN+WlqDplHUqmMiWWN9zbamfw+JVImBPDNqd
CYMs6EBsgYjvAPyRMrqRjRgujdM8UkpKA40wjIx7bGJWMbFNGX8NdnP5Sw04ST0wQUAsAypq/IVR
0ZZK7xzhBv+nE+5sII0DCNBFGxBXrjwZMJJ6AmYeC8Ob8GgmQg8rAYYXpWIJGTxoYDT2CnXdGkTF
JWS9SNveUQU5Cdn8Fd2fEhl1ClhGw9k1jqwmbOJcP3AeExWkEOBnYdUb/L+Lf7r8m4h678UZqLM7
pILwYg5AVeUTlqPulofuHthKzmRHY60PfQ3TqQqxQzChv81k44cRCqViMwb+9sgztRWEXaDlh6m8
yP7nlaqbY9XiQA+iFk+fnizg09IoIBt+h8f8wyj1jdtPx5CsQqjU9ckqOurgjR+6/DpDCMeUloP+
BsLeKc1TF9E6L9FQD7ibAVaYYzPCnd5LhXShH7Mz3a/RwpjnuOHQDD9BJLJ/1nY0SFyZWV2DOhaE
hix9BcoHutZAdpyBVyyo/fmhAl4vMyqjaRG+VTChdro7UkN035zQ+9u7MZnr4lF/21l0WrbxJJ06
WPcR8JwAbvaYbRY6T4WnjPqaLzJCc2IAfe4WA8FsqVKB4AbbuplKasSwDNzwzwxNdENTUjXdgR+L
WHOW8JV1RN+Kd30AWo8rnGpAastobwnIrYA6JcvlNWgqNYE4fvRXvn7laVt2hFV1uaonQdUYuCE7
w9/XZLV54A2+DdBbFpyzfuZUUscOF2Y9Vtwgec7bj8q2il9BmrBa3saQFr+AMVbNL5UkEMdA7KVk
v4BwYNLMJ6x8sP63ZqEdZMBpU623+TFKyO+e5cnVK7S4BW0vKoFjq3cQyC8szBxO8duY8gbNcM4A
96oRRnUXTmrD1o0luz2butuv1hEfxbhYHV7JuFvas0jOJF8w94xDtvkWfLDBjUOB6rQHc2qIqPiK
3z8SYNZRiOFykwl/yN0XsG0m6sw+RrJdSZykm1bOsfgTI8YKSQzqdQsPmmrRPChd9zpzHK3fVx96
9i7IBaLmTOLpHYj8QKs1r5EQZTFeCOfCTYm6qyCRIFBrptCMemtpzTJvxoCB7yQ6m/WLxqMdZG5E
lbnp13Vsh23vSyesJ6hufqYK0IBpGKPEWnnruKDASKA/EbV3ucKIHv3Owl0N7fusTB1y7pO0LfCI
MNnUgmrdPZBueZeXzYOxD/vEYxYDEeHjqsqy53UpUTsYeZ0/JLEawwvJdVsgJeIMtCmJDJ5cMWb1
C52oFNie8yuYH3twtTVIIGEKYd4BPkpD0cPjFzAs2/59Z+OS2QvYTmextQ8qsfil0Mu+WjxRB4fk
ULiS30JNRy3r8CjQvLjfvSGpVT2NU6stvD4Fq94LEig9zri9/axG4kwFs0XVAMPgOGbMnhwYPZF/
l9MFow0Alv8yx6krU1kw4sKDkn18M5WQmvD9l99Ci74aZVJJGdv6zaankokZUqXcD7UFp+8k/pnk
SE2asS/XGv+Gfg8UOtuM0RMtQF8P8oSX37dOQPuR8kcaR6k6/i2Lwy86be++7cQYvT/S/UpyDKSy
Le1rQRS/MpMaQd22GQz0KBlqsIJtD4s1btJ6nM7eoGZOgNfhzVSBVIu7166VxMAF0PbDZNLO5nIz
Ow6Fo9S5sd6KYh/aHBUGe3breNHArjN5LHl8Cxunq3prUk1uCFtrefqzNUye25SPx1WZ3O/p968d
g1Y+f8eucr1ouy65eH6MJWaDqWeR1mx97k/mWvsxp+3NfjVGJ+F0H2aQfnlBAg7R/CXheBgGM9xA
iDMAxcy5P2HHvCoN9Hp9OTgAjWm/7FvLJTK+Y/IECqbEy8kys4PPCYnSI0YegGDIhlhVW9NZnvpU
QWnm8jAus7W16ZiccRWSOQMpMBOkaInw6n4WB2bEMoIW1LHRtO5NShdhzgkvNJhO76Ks8zPdg/jq
VKSA0/EVy/yw88Km5CthVGWdMBBP/+rO8rQtzXaCJ2iK5G5kuTqAL0WkGx6P6MOv2msywL8L5nc3
1gGi27ytEVfvNq4e6M8wGibgVzo9vASvjX/zjxHTzBCyEBP9KGvGwUdUP9fZIVwNJuFc+Hk8iCDj
xdqIiYkui2Nbgi5ckIwB7fqIMhJaJCUOh7a1GK3GxFwl8jnDW61dLYxMQSDcUQSPqCer4V20pM/g
/ME/p6FFNxzqLQ3CzuFhSyD1fh2CZDskCnEbI9XwHkgH74dpxpN8u9NFTk6ZnZvdk1GaDIhm2d5M
ooebRGmXAb0Ta6bWErSiZI1BymWV7DwUmC4XXSPISY9KYIh2Zyn9j28lqM3kuUyv+5Xrja7c9jzj
uBRyeWlnWfHpI6ww1dYsio1LLcDdTArtlzyU43u928OPUeGZBhKT/pQnaKbr5gOMLjPTcWQYa68a
Y8taTJjk4TD3h4QluPP3LzUzejcs4Tgk3pgM8S49+enDrfq/p1fZBMwB5W1sBpoje+GW4ShKNsQa
3YFlA9vrcEU6tgnnRHfXmhna/oQ7gZxe46BYKQq148PqFQFb3Q1rCkSGMWcINKOLuT2/aTzD8ArQ
lvOUlvWlPI5bMlOoeEFAZ45tiOR19dsinpgwqry8g5WX1ad6zgMTttXezlTxsXnkaTlHR0Izewih
g2iqwz36JGHjuXJe+yAJ1mhelE8WHz/BoHOi7Cj2XwJ2Zm39tTx2leNVE9JsEBKDXtQ8FRiAuVM2
NEWEcaFTpSGkmJgscCorPgjiV/MT13h15DxhthOlC6hyWF2cOJmg2JnqO+cE8dSsBkfzPZIvgaQn
KTyUwDZNka7oKJcpHsGyxYeEuN+qh7QfNZEVRolltq5D/DH52XQjD9R+jTi1fqTlBRpmjFv4mt8j
2BZLBqcHAisdYvIr+257D7VcKy33N0X6ha3B1ThPHNvvCKxSa0wcx/vOCFh+qTmWYi483bdITvfx
2ziTZCxyHNayy0TETdjj3miadEPknTFsh29GlNX9f7vBltlm+MZWEqnberS18olL/XZK52okO2Xv
xFspvkoaWhNkz7SOYPnj7OWCftGcYPIOQVP5YAvQyggnzhroPH7jxr/SpNhT7ascmjfZi6LuYF1X
3EC9lJtU398AsdDhhtqKW8Cw7Scc90yJhkv+9Si+J+EiTlyly8yDX6KMZ9ZZbs6pgPLnTFT2fi9C
7+OUf4JkLmxk8fu88V1aORYmIA5EQR67PkAE9ZYgNpaz/BR4ub4TD21mkjAYsM+yTsgSUeynxgPq
bLh1U0gTjFVn77QJwh3ybwAj15UOzGgnX0QjXsUWXmaNnUzDHPLndvhEVRMD8ejCKOVNU6zZDlpe
+7jApdpPBoXIiDbK2bzRRSrUi0B51oPMWDvqRgEa9aw/Aqtmw7DNogl2aDIb00Np9zUcaXYCxQKu
Lpv13Itk2SXz731CCCkqaI5FiYa3okPw2eixYiNQywIgXpdM9RGERlZGbjSiC9F6nAMr6yD+xTLV
vcROsjZSXlDEpYytIdKvQiLWzhcp4mqf2Vh5o8YDC+UQrbn/U9Drzn3iDiTjKfW5oRkS6dQ3pU3u
Gxss6pR0Rom6wRm4xPzdMKZ0ry/3SnsrE8gUJWNvDFuN4foGubS1I+rNEs8gj70Bwt2eFRKjsGc+
IJt/chcGqR6NPatycS2z/SPrCoLLc2Da/q9oV6+3MQFM6PjoicCjmuRE67AhuUQL70y0XpaCfZpK
IAaXncFqlOON1oegmbNBMAaKqIBUGfGE9N+7dkrs5vCD7J9sIiL/RlR8g285ukeYkztGQ8Km/frg
gcgxPxygOrM2YwE4khKZoGmrVSFSqaawBOTbgSw1xd0fX9suuMYYaTQpbd/GpGAWL8wHZJQqFNQM
WDyQW353kHShOGjxxTZlewHabYioNdqFa+Aek6cOKnTsLYqwkGSjOB+rqIzgah3buyXewASSmmcB
S+YOW/UqWCdM8tmDzLR6sEydmhbSe120i6c4kEIR/Ldf/CjJseQi3tS7FzXTxcKtLkLQq9+prI6P
YZ3dOuVRGtBWMuOtkdpTH4lF0sNMjmuFtm7LjXnP9sFbjl0zKSjVYAjtCLm9anCkx5UmlCvBAjnB
lVMpE5BuyU4F82KH6CIBI09EiRCoYTv2fL7nGLFbjcKV2li6jXqj9465rsKFqv0q/DuekID848VM
ZNlPc5XS2tfJm+o6QO+eeHAmh5rUUBe45hs8cyV484Vyl5LvflznDzLy8C0xa2xu6Brz78ZpXsJK
YhVaNmq9SMM3KsbI5FLBSZgzCAmaq1CndUMJwB12bBpt7xnxTAZ7EHIr2d7ebTpVietS51ArEhJQ
5ry5VGBOM+rozK9oOewLOsjTGnZhoXpMLpM99yxe2SRVPqAi01bSKRIIPvSzbOS4dc9KePmhHwDl
1uKDLGMUV9g5DNtIP7ay45XaxgBIThZp7+Us9Tw1xIUjfQhYs9cS8uWvsWjHeAIpu13OEYQK5J5v
Q2n4IjBMVBBtKJiS5H+qg9/0AOklWC1rqpo/0UHI8FXi6/UGZORbhc9FXKi1QOTpQZ7LL35lq6Ae
tlbNoTtaa427fQzo0MP5mYb58HaIqt3seSGhr7KR76Uo3q6frYLJGgLjyDwc/E5eYXleVo5wFCZ+
ZZ85x+BhooLQ+Bwv3x9HeOLHLdsA9/MEWoLEC5BIy3tCzfxxQhYLlAsimH7azdRdyJ4q4fQK3HJ5
rWqHh0YwzuHjnTllleK8MKQ///Nlb2ZW0xIFR8hB7vrJ42OlVJ0CF1szAC+1+v9WgynaoMO9tGdn
QGG5cO+JL/jJYqymxZ2/VWcPpIyL4cKYu3VJUcF2SwJwVbL1H9rHuz1BXVXyDPmC67lu9WJJ3iot
nN+U/PSgn+8SXMPxnJxiwRo/h5QoFo4MDy4KPMS/80Ray/8B8dqEHtmRUOLWn2gLPSC+W0+xty/B
KbPSQTQykGxVgxFjdk4RupzGHJ0ef7UgfJrVLwYJWE062gp7yvVdiHWxu3GhtBngX5iCod5sYbY/
ZHmaurZddwHr2Y69UUdxpNifbUaRQ1UMC6nMQa1ctXs/XTE8i+bTbxig5FZxzeMlGvjFQVPWfKGu
nsUsMiFhsLmWSA5ALtef51prfW0xCTF/+bCrZPcWd7yl8FjOoVc8cOVfKoPrAdykLFdpMGI7yi/p
w6aHRsu8DUeoj6qKP+/Uz0xtiPH9YLlaiLZRTIuE5zIoxBQXnUbU79aWUmTv0loYIP82TB0BxcdG
HvYsP8Tgay9VfVa/+1cc75JfOD6WaEBaOk0PqAqwi1sU/CVUlhpwHitz6YgFiNb++OdYYqKEtnpB
jwTg3XKJVh7UQNZtmOzkd17MkJssMU93b97iY7ePVGHfrvpqmsD3wUWRsM0TLYkknJVfyh89erNN
rjaWlSzi6E1fkZuaLK4YwSKBjWZS0koW0jswzP4sE6MU1pTFeq76umlaMc3EQYoIYGnnXVhuDphb
q8KZjh8wfXPYW/YjTjtEUbLcR6r0GgujouWxZdJiBAnJSY7JpLRI416VK61AU1Ka64VHm3AJWSGe
UvSIZTHJoqzhuJghohCGoDYoAqlG4Mnn8MGnYUDbwUM/0KfbaQjX+rh/LpK51opm9ewZp87G2P0F
UCk5deJ4vf5Rz1Eg+I15rca1IIDDKU6wxZTLz+YwfYl4on3mIestSZPRXCiCHsTpLBi7imKwISbF
8sw8lm/Meb56CMxYo1l1Q0Klr/izWI5cr/ZONYZEAdysPwY/crpwUC+TTkekjKRQXR0jHOWT67Bs
L9QROl8I0jcayvNZfzVVFTYVMwoCaoG0oYP/B28ZDSS5rYx8GRtAIFQvwKL1xe6lj9rDOF68mpOp
XCqYeIbsC09ltN91STFwQUtVpYSjhRjnZWzsg1aKKlNR4y+8jQfI/SEBTZ6SvRVJs+1xAe9HSOXK
co97Zfjq9yokAupVpAcf1H6/fsDfl2hloSLbmAFRUfnXR92DCSpnKuQ9O4FDECNWQIn4wVNgoMb6
anY7aAbB9a5Z9HlvdyDMOUmhpEkFG/snZ53CdPVgTY61Ma2MnWiPc+S2hR5DsOCc8UDc0oyglpKG
qViS3zmqlVQn4iKQ2+cEgH+lmqzaOArKI1rABHjRAf45VttqQd2uJQcPwz0prpWh1Sd1JAQ6fFTx
HPvgYiw2rrsSouLhalLL+VXFri+IldTZZAfh6PvwEDSBTRsMs2YwbnED1Cwce6xPBfmRqBLc0I8M
Cm1P1uBBq4PVw1KG+2zDqCcnvnXQj//ZjCciANoPZT7IS865tDA2dJ/LJFvjyB4Xdtaor5ra6Day
A2O9xAAAZ9Z6/CNS58pLa/indpklrgDo2vSZ8RdwQ0Lr+YKCpM9cSn1LD4g7ZHq3LDjMIeOtdHK0
KjIoL+2USvKaJZGi2w1XwKpyedI4C7d1KJHW+4OQ9jSyRbl+sUjIrZRKpSYs7tkATS1uLcEolAWh
8jU7MJ70e/r8ojQX5vdN27fyLHiVcizsQ7ka30YjLK+d6Qfo5Kzl9imkISkKjBuhDlzL2Sr65bb8
nBPF5/NpdwSIMWAjSUkwJKluvcOVmZtkBBS1v6vpAwfXSEj+hVJPCJ7nqrs35dQ48Uq6QhXWvDcR
jQgA+HAnLfb7OsyPVE8mRYOH2l/PN6/LClUUL4t1tmKQ6YVjsRLQl+XvCWD6mRPmOaLR7RsKipn4
ZizSlA8IVqpM3rK06T+bVFHmqysj77dFMkro7gjYUZ+DLwIASy8IsYNSC7ltj49CRi1bQztbIQDM
h7qzqIGz4tFSrTlBG7iBhbJryJBSpdYfn5Kqy85oYafEoL81LfInDeqysB6RBBNSmgPDqWhr3kIO
5KxP31oGgufGR/5tAteibOjWdWIZ65m1RToy1JSWaZV5EsPDJ0cujfXP3oQ4BuFqLlYojG9DRRaJ
r8lReuDeISAYvNeCje0FQxAAYnujj7kKW2Y/QPv3KU84J9rCAMLasnOxd+1wzIiPkNOT3noTGY+x
7P0Z5gq6O27dEMJmfj3X0bj0i7v8ZynmBEIBpv1NpnPF+SMe9GCgYouVu+KwRZlJ2wkJD8azKzuh
8XZ2ULw9lHcRsYZK/MJq6ygUN7UarwGwlmwy/Qso+iriAnV6NQRAzQBxzpecMaZgU8AdL/7YKDxC
yPxCUcajM2qrQZ7Mpz3yNvX5BS8pHyaihvOGjxj12bIqF+df4XFPcOZWJhiJ0JIKlKS10bJF9vjG
nK3v18Ny0O3+mP4gfofScy/6hve6+w/6DHSrfZ4oWfM3gFcw1thmkphwOOlxuh1KfKjAH4MUJlyg
NqPNn2fwuejYVKh1Tu9dOZ7oSuay8pHCKIqx+BPBQ1hrNgCnUz0QtFRlcZ5dDQ5VyQJqyBW49/pe
hQudHfdJ8abvwC7EHL7gvIpac8vpFzrAgICcU8eVWwy9heJFDypETg4F8thaEnJI41R6ZMHQMzkP
+SJVLZwf3IDEqXcY4rmftRg0/A8JDco2kRppIvDiRr+Q/iU/D3GjQeSUyFTA9QpK5UYkTUsWpJam
jgv/WPXRyF1IWO8AbFWB8a5yxhbsMD9x2Q+OdtJTo7Moajjg1YCjbvD5OJKGG285bS0rntXBd7ca
kx+BNse6Gd6nN6sTnyeFNcy0xzSUli+swelMpRdmQ8BnN39t3AXyTpJyD2tHxu+c4WkpxLWW2OBF
qDu9u6EVujb8bh1JmFiKsBSMLKmGWdjaOcYqT04cy4WBdB0jR4S5ygKKpY1B0UzG8mbl3KP1EVZx
5IyxSMprtP0nzqQ4w1vl2RbDPzb8MRT8CiPiI7FiaOyLOe77YMP3ZB22XlP97sL0Y/75C7RUI53D
713V4Yx0qS1HhFLhmjuXP8mWhYxzTchke2YDGQaCiXlE2Qd0Ryv6AvFy6lQIuiACLiXk1KG3XJ68
evBRtmksqTN598/V7ob1iLkcoZOiu7E+umas+/BEFxlmuPWknsRt87Kr7eEyYORZU6J4hlvggbzk
a92NOJObezJEIM5ljEMabCVJPuzSYzibcHrw+X8s39H2tfMG8dHFo5UaPV1DS1kxWwgk4ZC/yLHe
8Aq8aGdU+xc8HbuiPM8VSan3rzJEYQaYcz+pJf3DmYAwYyVeMHD5XpWlQ5jaUt7ot5x3vEWQuZlc
ZDG0EyDVLe2OgGJkJZ4H10y01/EqK2E0PxerMfxuu02zh+J2VdHk+t8GHto8E2dVCjSCPyqBEk3U
8IrflqnFvxJzqXOmvNryT1Cd/9LcT2rVo+xNmX/U6kg0leclSKXFPJYKMxTZgySMbuT1xEF+8H51
aW22gO4YZHOe+Ab3IRVfgPn0Jc2z7M7mXnBwrYrcDVRlgmXk5RGeBrddDy/lPWruEq/DrPasTo/c
+ARrEZ+zIFnI1AHv7EvqpelpMkfW1RtabRUDfG2biiwes9LBYQDJzOphD0pGJbj7wg5XAHxVTtEI
CwHeA5tXTm5kxD/vcdkZNAJ2MdibgzpgF5i/4Sp5t8JLFnVaq5jE9X2Co5e4l270D4D1gRIznuiI
iWYAOG2YPW3C0OpMqSvI+xzuq7hCb1Bvokswj4qUxcAmtr0A3WtkGFJUJlg75ANHr65+0ZdKNn2O
5Q1tIw4oQhCPwNjggJzguqLbYVLLYKH48hbjRriPZUY6g//atqXeMLki0ZzkmTwvHQOItbv1MCIn
4BrHor1zGK/vDmd20M9GJ/IWjQo3SHHPKF0xJSuXHp4IKsGgVoBX7StLKsnaLM5GWhwgwpw6HgOB
wsBQ85QV2kVHL6cArtzELJX0V8PAdlsZeCA/r48SyQm/QAaZjxjrKPZfIB42bvzDD6pr9/zSCDJ8
9TX6rRwez9vIcoWkpBwJq24zLlmxP39l1ZPaR5AVEAw4J+jonrF0+iZQhNjyxZRmgdgssgXNPyrP
u4XzspeGXXzLVBoc+8rxjFqHHSh6FPXzArbEJUethwetwQThHCxro81j0D8AaiFv8ddzrhY0FNb5
EsXxe0/o0urPrcUCk6C8EzXCvGmhM45DTWmgAzz4fo+7tH6G2U3NqK4rbj94Av/P7gBq95i7XkkD
G6RBFkjmTR2MZ+8VbUKvITRSSMOfNecJXGV4qKNqP+wrX+uKF1vVQMYzNWqMj4U9dbVpmv7qyfWI
nh8+ntbnkeacdl2TMxf6mfDSmUR4GDqRr/+dPPdgiNZmjH2AwvBZ/OT6UEpUkCvokjWO0Jsk/AD+
wd2sSvUe8u2OKkWmXg+qdv7etK3Zzzl9h3sV4CpRe4A3p1qxD5BfqkQGQgQa4w4OzVEU+diMkWq6
rg/gKKkwKvdWXwFJlGTCnRY26f0uEp1wZdl6OSUqSsJzALwGjcXfvOK7cU+a1UaifvQWZV45DN1l
iwrHC7tGmVorsFBljr7PdJYgb4eM0X1fA50RELnR/OGLXh980zFCobpb4kQSdKVR6l6GwEMtZZwg
g3VI5J3/KApsDki0oiohND40lRJhY5ACf8mGIu8tySTl9r+0Q7WKUnuIaSRrAEyok30HOSuDNcmg
PEqB01KnRfZet+OO+d5c6ERzJNREY6V+LGSMMs//WhOK87CkVByM1ulssXB/uQJd/LIL/LlT2iD9
QoLPw5b1jpEgxBzK2jcw3vHTUjnwv0aCxohookjezLJyEeS+6B7LJ8MacKTGe4sxnl7oI8f2gp7n
hVCBANxLOdzMguJJAKn6cG8CywM+T3uS85nu0H8f1MZefex7cz7d3ohla7Iwg07jMyLJuMorjaQm
zfeRb7Y//vtEN9uDPC0EeiLlxeL4kKgVDwD/Ipbe50xdFBDv7qVHRjTA0aJJAE94EUdAKboertei
Elc3NXUJFWTev0k4BIRFw+gOMMVkuXCIfBdmt/oqW++eokYNgH+532h1YnbY5bq0PaRYRTswXL/V
W/+FqgA1Bi+opNcmZKHuM8rDVOa0eGBXgSeco8OIJPlSFUJvTWfIRRqxEXtReNB+elt3oQPggVft
ps8wySJFRrUpcSYku4LaMCkJ+xQ+UeuMH1IZdaI9ffRRgRyXqTw5HeVzBGLGm3j9MevT3XS5ns09
lkGqP8fkjZA4QLuWmL1rTHlh39Y1IR5z8C0TOOsGL7EV/jgVr+0rfciNU6l3sjhMEhrE3RFxNeEs
Cx2wWB0+/jjdGzwR2q4xfdBdfrjFAepIatgEWbnPqZrficwgHntwZY8Af2PcA8AQb78+XBoLnRor
GelcwWmerFXsVuVEk14DQ6kYDVPQwwe1P79eESFE6ceTLFhJ4PpZe4gSmdM7xHl7pb2ulNKRLwjr
DD/GGYcgzoXAdcMQ3xQzuA90rrNEvqhoLiLPgkttJxVK7gMCcd0lCYuRJmMb3ysybB4gXnL7CeID
WyawHfoSzfboA1jxGvI3cb0dJikvo/u2LFs5vmOT2vZee0NeNwChfledD66HD8WS0bwSEWVsckXG
5cDEGXmrraBTOPKeH+scqw36fD26oMu7ZFfSJwphJA2C+qeYmnuD3dYwqJy7SstXvFHawnzmWeo/
ROk6LfSaBXFQ73dhM+B7bWyVjxUaCYL7Lzed26HMN+OnBosPl/dYIlAjXL7W7i0Dby4O9feJXDn+
hcLMwV9iCIWh53ejcnARWGxT3cON6mJ2g8HpdUkrmNJtLntNiIuPcs3gdG7MfUfE++kcc5WueR8o
Bmnn5OyWO8dWUx7wzIcCxUOfwOMwBYPQfpnZ0hTJnfojx+vRuP63jmw6140q2nrX5slhhz21oibT
8if1pdCacPttjPMk1AaE5YFrioN+opvseaRXJE5nAA/+za1l9ibxjKmKUKMw3G87OMUOjkNfTlAk
B8qzXq9+zYeaDKTnC5Xt+qwmfOgfnbcWnHggb35Yeb1XIw9F+vkMwUcWkaWzvd4a6aUoogvFVOW2
r4zopiixpaf5YoCKNSRo0xuHZW6QW1M145wlovVxPIpQfaT2HEi0lLiJB/oFwOezWpPBgBbfw5+k
xG/+IA53vq2AK3rVZCoD/6FxpXxt4/EnlU5dUVwor6i6ZDk5dwUtxXWDjuxK5hye+XDLc4q7GSDn
fubAKspOCmc4UzrCCLDlXeSjm83I17UqUGffbpMTQZ9klTNOxWeYofIgGCp8tyiz63QmwKnteCAU
r2jZG78Rto8eSVrGj8r8OvLJRmogOdiPb8C7shibZPhl9VuI8U9cthumHwwxA3q02xWC3nMvEdxC
6Jxg83CdNChS54cOdF0pqu18unB4j0iB690lfpw0y1KvfTbDOSSYDu45R5YK/4lqGsmxqjuu3bCs
rakSAndEZ0dvZwaBNAd2paQzEGVqyUNUpBYBENtF3MrPkjvmV84jSJr3FIyIOUtxyp6IaZWsmCYK
ljF4mP+Kqetq3rt7EZu9BWi7l7Eo3n43WAqi8vh0DmKWfTgZzri4CR0o1UphDAWLAZlRgpFS6qi3
GVzHyFZoUp+aJJGtIwUSA/QZGfX60wlvIOOaXHjNID6aaRb/Y4GA5v6m+VWQXm8KE74W0R81ey4t
8bFfhsqBNVk3uib3x8LHRb/g9VOV6XllfPuI16DwSaPiwFySrFdAoBhmoD40+Ly25fjXoVfXb5+l
WfA5+WxhG90beGPnVOMCT3Ot+tehqUqWS4RblmNvdnVSfxQhMChnAdFfdM3IwOHfpWpDltDWlk/5
6dn9ryfF1yKEsM3zS803/tACxdsazHGEWWHW14hP9uEKETjfT5YAf+ZVOpmB7vV/smTa5wmgJo9W
nTDS7gN6YVYCLqCSXIhtV6Ft0QvYotI/UB8NK6aiAlJFYPNlm7otm+dOQSzRdAn5JtPjxCzeb3fz
8CRtaLi93WtSd1L80YiDu8QS3Chp4XpmzP0SrOc5ir/kdVAQlSuec/BPb6+5MB7BCrBFFnsN+jFB
O3L3o58GUaZhPblJZDHcAZfosd4viZ14BrjOWklDLfAd1I4/bJnPShqPVnMdcAKhiRGRPTqL7pew
DdVl2/mFSoVmwMvHRxKHMEvfhv+HHb/jPlGy47w3Yj7gzWgjLMAfpclwh7nmlyAk7uGOcdVD4eTj
CJFCaaTukGFDLg2Mz48/PDOYVSU502RsohZ1zn2w48Az6kGk82k9nrIxg+Fy5jrPgtn/Dr4rrWl3
pKPXFuVwgRcncDasDu3xeP9tihC+8t0cbxhpi+kTwRvBDrHxyjVkKgViMJzEc80R+Y3Xg8TYcQlJ
RSBcOI1A7flAouK+sYTQ/rx60Iufo2XCHCFirFkROFrd82Ar5q8HcMuj9AKbRZ/qm5KhbyG8lzoR
c6ytPa+lZHC1QQXNBCFgg5ab7HF/wdBDP/adG1IrRRiGNAW3KQM05pjTtoCIXIzZuXWLqmqvVQvL
rKGChPj59q/ojuanpQlJN2KXow+ESy7GwSyfoXN/msmRegMNMmtpKPcYLqLqQw8f2005cvOJTJ/a
zY+6Tk9CS1/BBQO4w8Ac77YmHyMRETnwc6jmRHYwhtG1URClDzYx68YUCdZgPqnuxQ8YmeR1pOEV
m5xvCqBUm8avLJD4XiCCgrsQIhIXu5JJDaUmbKdXpzM/SiXun3MLLPfJVivZu9Brm9B2b38pj1/9
HJdIQLeKjlirWjLDtTlC9undeIdy30Wob/FemcBfKIhEZ/XGKACSg7SjqkoU9qLZtFFqyncyQAo9
BCjrX+o7EPsp3Z0mrkGtByO7pLV44B8yolVEB9wiInjdV5ssDCIt+e3QeIBgoEymc4+m1pP1uUI4
QzFX+tMy+9hYtsMydz8aF7LDSyL0YP7I6uuSef1ymkEuUF442s3+7sWe239sNj1ieL9RpuJNfBme
U3bE8l1M79057yVJsBu1pwZxKcJO+uaX7v9oWao/Zno7CqWBzxdGRZs9Sn04xQ9ou3xeTuIoaGZi
x+IUVSfMH2VwZxzV50ECzHgPcOgLDFJO1e7YN8EY/jyX9lMTd9I9m6GnsHwdxiCYtfG4cd/xnFTU
GN9NwEHUSlB5B2DAN9JmAQYPxmFJKCv8pCVz8k4AoY90wMVZ7gQFDsi8/h56lRKwMYIOYVh7E3qQ
4Cu4pTrTH/t9oHyGzj3gqnlkJKECRckH7nE1CUTT5p6hN0fvOpbHLp80jTDqPlOZEaSesOsmkZ7L
8k0oBYLb2/RzDl2AN8ID09H+man32fr1eEAB8/scPSzi+g5A2LsJ0l1wynTJNRi9c5rtWXsBNAm4
v1NTq76i20DFZkADYo/p0YYKSGElTPocTq6QqMEenXCyWaOvIGAKorgF5Gte8pe2qicODR2O9We5
0ar5v1CHSrSI0mkWvVzzqVN4bj4RdNd36ibzzkwwnHw7a70dxrGGL6W5IpbANjMeu2VNKgAZKok/
HN58lTcOtPnSQdQMgFvkITlWJYbzKnwfvUaz/HRyyuQL+bF44ILiA/McvKv/fgRPru4MwXmJ8Ett
sNb2n4n/adlsfPMjEOUjzhvhHgEUigHKYA2YnvInaCHLUAFx3anAeIg9KPiNjmWFRsBcDv0s6I2e
X/YzPEPkUYejyeO57f4rXp64DlZlYVnVaO2duisGRlKMuMWgfJmayZ+ds+KEykPK2w0cmoAjrx4m
FGd9wcblIMR5B04ASMbMd63nkc0L1GlCe7TP9fkNnsov0XeaAhg9c3iL3h03rzXmLA/5aiVZo8MQ
vOjCt7Cuip4V3p9YUgVSrXHctJumIg6ihYbv6Qd1pnWUpVeLK4qZ9I0cjFQOuVY/MX4mSTrsELtx
QBgkvm8lKBaSxx06Xkyr7KZwIvhmEMqD5s5eEZhJGm2yqNR/Qoo25bCTuA90FbT5opx5kszbtVHx
cnfQso0cmf4qlK6KYE/3nUKmDvpwMRRfvjNwboM+yR58QggNW/taH7nYy+8OiS1UQALPkwqPejAn
J6H6DvQsR8q8b8nxacXBc3+N4DADtkcJUxyo+zfF4l5+XYoxUAUbQ5esuUmDW9Mm1bHlFcCiV4f6
qxZBvvnXR2c2115T791vwISewqwPgRLW3+onZzogktJRuKs392N/qr+XBeI93rPcB+eEIxx26Rc3
96WxN+SL4fNWLiYdeMzCbFsZ5CpBD0fX7KarJ+F3CoGJHQfHnkgZlTkKaHMLX+248MxoOknGFHtc
1/kn1GD+FF8vsRn2yyenHIr/AtoBRTGGRYpqOmYQc8ghc44Q3EMAT9FnSWgS6Km3igpZyFZ9sdd9
lyCz+4oOJYgrS0jjvtejqlY8S3TuiHejP+y1kCUf0LiWcZTMbM6Al82BpaR6SYAW4QIGkD9MIBfH
ycjTNpxe8DZq0ODa7Qm0v/8Kb1jLTi1HzOzIRDuBx4niO7yRdgtwYJ/Y2+npAe6qCmuEUEpNzH8r
wJ3wrRjEC9xicoqqgrP5re4fmXb2JHGtzZyLnNmGyz9PCKqeLKdkzLwW4j9/LM1Wsdc98o8Us+9A
OOQlTLNxC6Kq1Jn+ECbXgfoYRbKxMXaWmNas4oswKXuSvPyW6t5ny3Q8DVLPZiTQUv4vyPHv8RLU
8/eJncTQylf7xii6zvUJv4AE2CANzmOYztC3/txKs4N5cOtP2rNrsIpCOAjCg2Q6zSJ61robrbqa
J9aS4ZwMm35wZxC+sooLUHmSFa3jtRsaxcZB9hffg+aR7p6e11WWUS0IIY+QfpCPgOwOKVKm0rDy
+lpiZDLAjAliT9wKdcMbiq1bV2H6kAZDBxgdzyQxr19W/V1Jeqbk0xKMi6jnm37w2XhT98KJackj
RcDhXd4rKdFBjktmT032nEL/YLo4QaWf1cLEkBn6w6b07hWrvPvXwZPiAcRIHWr/2qjhUkY9QlgN
6un780S89tFMlSxsavT3Cxo+Gy8ZP6DCQe1du2rssGT+1TjVr7COPXVTCU78Dck0Bk8GtlzecfLd
cblip/jDsI10FaVD5cPXT7UXz9zJOhTxd2Arp7HOW7KfOGy58MvmcvsUFLvsSp/tm2rwieDNu+Da
VBo1hwetovGN4/6dAAdBfA9apPau3w8jeLCEj5LFbq7yAeW4TB2RH9Gt7/9FE6aQduh3Yh3PFsCY
3XmmnHT40gYGo0yJ1COVl508ITtV9WVPiP2sVEo83ZmVvXdzBpVPrAycHrwSwtRxuSIxOoTIE+VA
eQbUTbkWKjwTOaIv0KsTT6Vq8jUrqQg8au4v0lXrmW4hsPJlfPxLydWDY5GIxjSsxJG/SDHIKxAY
XLj5wroD5bnZTtyvh0devh+XnDMIYvevVFnDVt+cbM5qgV+aOMmrHLmmf+j/WpLMOGg9VX1jbwpK
oj9xwNKMCAsWyYXTm0ifu+LFHF7VPrxdDFe+1asgPj9Pf+JH0ToeOEG/XQ1IMme4QbNaQHMuGyGU
ydCPa9we46OYYFTtX6zftgJEifKeaEsUYooJPxqNvPLB4p+VUQqe8GPgpTps1cdb1frzobVf1VpM
zEta94QQOKHZbQ+4FCza48kQKx3mDyrUEbxvSxJ0xFhPWLqKWz6+yLGSvvDHmx1x6ASyDkeS+2Nu
JXUc+UnM4YkFsP7weQf+R7ONJjXnMpStaX6QXrijbAd/Jm9axdU3goXCQo0OQjtbwE+6Vck6uObW
AdTrzxVoRYG9hCy3cgO4FLLmD4RP46PZkTwiUtxoYsH/DsbLrRVppY0nD7xeVvMC3O56fvHxFJM3
mTUBH7pCMfuyKKIyMdZW1ud9uMFCP5mJOwsBGu1CIwlz+1MPK22O4Ec4bZ/In30rAXqBbxvX3Q9l
a/5g87ipR2vOCFBrhOJ79r0WQu1MC0ZXCY4oyfU4MEgtIyQ5gZTmMbqD5GcGnoM21+gmrTek7ls7
p9n9x7k3pU8pZCg9ANyTBgToPWRBgkXj6vPvADExO3otSTrF26IDggObhVfew1XLFkmhnhNq5N2i
8LfEtEWZkAOwDG2PJeQMKGPxd31Ofs07DVU/PSVcseUatf5UWVft4i4605IXsowo5hnezh+QTmZP
qwH90eIuWItiLLZ91FM3GJtXktA1Gu5PYYNqehqnjnO8UnGi0xu+tmfsgEGGJPkCdB4Ku2gv0TjL
YRG6/Y96KByf2MwJ6zMjbUJlpIymICubZF6FIQ9bJptWUkFhkVqWjgqmpBQkvkb9dpWYclD0HcM/
MmGQ/yWkAvAoFZ6bSXRCxXFv9mJyuYxlMeDe8yx9E1HkOfjtDGVyC2qu0K9pLAeomZFt63PFX8Go
LTrBND1/AlCHyPLRMRVhIXbgZoccehs+/4f05lmw8nzushyvq5MsldLeuJkp8+UK8UuC3rzSi6Jk
bbxdk/Yh7FGaFFj/rftkp7Zhdbtp/f6HLJnJyBk19/u6sjAxKZKNFfYmh79aZ4/GLNjmwT9P+v/k
q0E7ag5sQ9Vvx2RF7zZnsnd4GCRxonk2d3pAywy+uM2PdRM7ULGRCfuBd+LQE9utzuTIEsAPH7wm
YHruuQqZh98nslEzzqWmdVa2tQc2uxCd/7fMXTB1lDfkK8CAFArcGZ7DCe6C43oJU2IxlYO/S5vC
pdsPx85SnnFv01c+ZbvA4FELS3x5O+8twZ1tbXpnaYwEAV1INpuY3GoYksSUHAfB3J+cE3amBQMp
NQnppIHP+YHybjVEcrZvowvyBQzN7/bSsFam+MSvpNeWsWSpa++//GPK1xS1jUva7Wd+DhP6qED1
yyu/fFkyJztvDroRl6Hx3rO5fbAT6TEgeJQQnl38Wu3usc8IJsmYxnyMPcot81QbZnIfNo8cCMAH
jmRwzrz4zS65QAZuv+f7L8HvsyOebxRnvc6NMk2CBrwoC+p8GmoVr8JX0R0Y2ok5aOW3ZQyOCuq/
VDbZ2Q6UqHLwe4q6isjJPTB1BOIpQ1+dWNw1u5mF31x4CYjO2zQIiIWJzjPSbnGTPAsvigzkxxZE
18KU3HPNRoYNl2Wt0jOpQMIKp7JUd5inv3mADd5KYnDKTKVQupNdiWTQ53iUfnLFDaLxHDsUR5HP
K3XgPKN6ls1ayugORYlbX0eYKxdeRRSJXy9LkJYujOxf2he1/GIHrSyj5zsWuUYEapkoG9oiObWM
XlvFFgtjr6LDG3aGzRKMMGjkm7bRF4TicHVTTQ2kOXzC0k0QvZAlpQZ1cjP28EMkyza8jEjJRp1m
csgJE+mc43kYQedul0kn6/gSBRfLpJUiWlVby4sAi0SaBQPFgWxKbG9+v/pRAhfiLlS1aWw5c1h7
l2U7+AozDeEI3sOHcgRr3hYq1OOVLPH6SOkkU4q4hmBXk0sZStxwks9I/z4PoqRl8sFi18uHDq7I
Xpsngwyy7QRA3jkAxDEzT6HkUZlXemAlzA1XWfxLJE8isq/6l9HBVxAYE9utiRfIrmazVCGIKxXV
lIjSVzaV0bOLY+fR54ccjMJWUwwUucRrzOH4l+A5FR5WQAQYHxPyEWAyqWjcjXnPjEaJML8+Loy3
SIlaVWBBFy5cSIrWpk4mP7nEyDN/b/WiLegHFb44OVhidNWx4VrYZZyfSM0D1X+osTMrwYFxUT8R
Sf04MP+JGqwAoKIkQhb2atlKk6p26WDrFkkpTqNFIqWJyeTyYPrJgEFVR0LRk0d5RwYSEsDuUzUK
F5qJUq2dYl5XkYCA7mu8FTjTuolPRfbAC8hvK3E0cZvs22wZAXljeRzy+U1U6FbT5651HzJPhHCL
QZObUp4VgmkALngNJ69cnH4ciJCa7ZOicY75PmS5yNjGiyEwzcgACc0fdRUxdsQcHLq0WVtq1aJs
FuNAJzo+/DYiZi5JSB3h7q0oal5khMoxHH8Q6tjydKD1uT/9t79tAG6BgQbflQjylLPokP/0usTY
naOUIMRqg8WLSQIQZCxf/Sm/CoEoQidAm1IM8TYeQ8OvTJY4F7EoU/9cKIocTspTz79WKHE1ZUhO
E2zB7ztJw8vCL+ELfyjvGRHjOnbj7QMyVgam44IEbVNvGoffhsTmD0rtBsiDXp+ozy8r3yeJXsSj
+awmAuxJTy125LPf/D4Q5dcC4WrEsyB8uZXClElCAWijS6Pjeo9Rdv0icNKa4+wtWxTKgPdPZJao
wDs3EPVUowfae3KIY6fpQfF80ojVmKUq1oTepHek5LHS0MboKNKAHKSc9Ot0XEFb0MFftBeUPHCT
wbVRgTm0AV+hiGEvqOuozGKvcVQNi9XJYS2Nak7wZamJf+Y4eWmB2yk5gWZxboxik5tPqBZLvpGE
r6OXeMBBPWKmOsgoYBrZrVmib821vI+9Xbc1WRLurWhF33EjTrrgWuMqx1a6XT/sHPxKfTguEF3D
eiE4MVgppynv1FH6Y4cDFCNhKfahgWsbDW826vpj/F1xkOqwLG5ioNcKrUasuxRjlBZvHKuw9sEP
0RB5mYABT58vvwgT26JJrCFvImbiEkrQJUUJJoMxymhRqLAgBN3Uvs/k+gY5FmfU0TsPqtMHhlVC
CoJ7ZsjtENbfKegAdVA5T3yxkFQ1lnzwT6BiLFxMBd/6uFocc4YAUaU+iRMKPs7ThTqLh2fJn7ym
JTLl8otXh9cqK8Cd7PvDgPpVFTYcxGAWJTnUsmCob5HVbMvJXp11NjXPwWzxC+NtnpW/Hp4c0NEo
+4m+lGLe3NH2yjEpffKNLkxyea5ojndHa01k6xAwv9orWIJJ9DKKDKmnujQsvaVzlSrHLNgmxFNy
Q6XtOLwXrrWKFOVCkCLkHnwdhcAviLKDHvGN8351znk7AKXFixl7Is0RMzFu+Y1PFigwOUle2UIz
4HWSj49GUQXgs9JqIjcEmMmP4nkPv0RXgc6txo9rrPjYTPzxBFKQJyTkcJ09Nb56/5/pO77sfHuJ
iHkN4bOF90QDZ3ar4XUnmH+oIvu2Prd/252bhXcaa2PkaI+DUhfrSouZMhUk4bfoBCYTD7Z0Vum/
upoTzT3dCb8F4B8MXZpQU4miS4SHOA99oH9ZTCF4mPjwThRgKqmhfGAMmoXR8e1gYZPyOe54D6rI
FX8i/vQjQHnavX0sSbqVxOxk9mqqd13WNCEdsZkzyjTvX/2Xt9+rRhX3LB0WW607vhLhBaGC8JE5
lGcnODScOwMMCStPZC7Yagp7JB3YOdKPDyd/jZL2XwtXCRby4my/iANWhEJtRbHI2fzfgn23POmq
mVNnRBqylr3wAgvMwOEt4qDklfv3mmqRhto25Abg7g2M0hrKeGLv3LXAqFSTnsC5cwKKrs1GCG4i
iMaWM0XtdV6SXbksu2zZLmYhuqDxD/noOghU0fC8hKI8WKAK15WD8VW49o+GOL5k7AMXuGKTStb0
gCDqNUenigZA5bXJVn/iTQQWQItOkmW0AcRlbn1MLsuBHme66yH2UidmNn41tRDeY1NYy54k52OU
Zk5mlA/BmS3ooq/l1SNSUCIo4FY2xitwyaSR+mP7kpuM+noNknP0L9IgHLvTR8lIMq4znVG6gJL1
EuH7IVkwY9PMFNf8j0eLQSiCIGtSO1BuRJQvpNfBhFoHmzEc0ZQ2+LmZsSQ2VZUrfe7Y6XDMLf2v
2LJwAvCzj1CBfo+t6U0IuZS5gEbV6+YkehTGix016lOquw/8O0kvbx9ns3HT+vVqsfrxY/UGM3gc
pB8LF3yrE/PNiWosFUErKiJNEOH+0/AqtIR6fidpvOG9Zmh18w8z5k11U5nvjoMeCsvsz+8Suub8
I2byBXQkJJo5PPGu/+QzBVFvjlJmcOwICSTj+8yqMYo5HYMbsKEQBl81+26cLk/ntli2dgM77y5j
I/zgF/yt1rEL6pt7dHd+KPre7Pw+kwBRM+1ChS2TykuADrJhc8tVItqkCNVNb/Xzws26g12CS4m0
Bwucf0rVbCP7k0d8llY7iTlJTEN3MACzZ18AT9CHzQFV6nvqf6mygn92E7GIHXmHJgHJcaQoknuK
xtwNT5w4ANnGtiGkPUT5fnsiYlKDz11llY8SqD2VC1+cRgMd8Os6uk36nzTUmmbxOomYOYtOx3ah
59HdXKOFfss09wtdoiwIOc1eYsu15O8HYlI62QNidEL7BrKFrO5v0S0asjnkWr7kh+TTPO1WWpjB
CI/q8c+COVvYVGifsLICiu5mJLbvXcWcT5T388CULzZyURbhBXluzvyKspqZZ4w9wr9zkFtdGQGh
XQhfLs88iLeD4PIH3JP9mJxv43HUzaFBmIYfyz4aIGrXqelEnh/rLiff8nHVp49PRRFL+tSkgrsq
zFRzy7XqgjIYttEwSvUBAn/cc+lLTIYpGKYRKZUFfSQzHcU3GtiJcEcdu2jW4IV38BBoGmiDVJEt
buvsabd5M2WprRocGEWOI6XJqIzIts2hLkXdTOBU4NcnSjOekjUhyAwfclks55t0ECRFnghOSaVt
Vc3mQPJ29dh3hF9tTLiES0XxSuPya2oaa1mVXEPWusMCNcdEMuObn2kJueCsOkeD8qIEW9zo3TFV
uanqIdXiMxHplHmNeDzthzd+fJ+eoT14lVMZNdqiNCFrjNfN+R29M3xkqffmIrNurwiz28Wx4/qA
QACUoHa7h6qf/Mt7agLn30lBSR+QEL/OQzM7w604/OBkvas7dnpmWlOfF+TBwMuz4UczIk5muk+s
gu9aPC+i5LRUTExUS16hjrgoZzPEs8r27TNZf4/rNll1W5tdipTB3Gz3OxOfMXOXBgGRPvSHP3JW
W+f6Sf6DK3n0eZsiUiV17HuvADgHD5xPftvoBIDsu/MgPm8gm83gOnjW2huf8phHLNJ3CTR26CDV
qwvJjWdoXsKpaCzrRepAhrpxesmXJqfgJgBbriH67Rn8Yd1Qr8YdYDcdh4WY1p3mzoqBaSZmmIA0
HFupRvgTjg5KEdECtBjiwdrmOD3mn53TGXRBOADEpiWBYQLRcE0ilxY4cmyd3ZbVUvhCkSk2PZbP
jbDZQxqRaT9dp1xezo38iYWlRgoLwXlUpa/BkzyH3Ur9sf5XG4gIWbyvUqXhFkrPGtO7qhjkzhcD
eKif6D4LgDPH1qBqdyhS/de0sq0l9s1xX2h9vJviYxWezih73EAZ7XVGi/J8rTmJ+wf1i1KRAsRU
ZC1V7kRLfOvhye6CkBwYag+ln/qB+W6WspBcGxAn59DL4SPUBBIz2HpO7B4VLPKxmg9gahej/1gi
NsQKILn7SWM1Y/4tzG1deoHtUZrcDaha0a9iMTgTI43ifxVyZ2uAVLb6NnvGaezzLN9HLAy9H8f8
94rME99KBG5nt7iQOeJdwqH4yGw5C7FHArO7/p9yV3NCAm396/Y+7vIo+UFlzZ3suSEy7z1bnWIm
JcIbWSljxirAOMT6lUzerMDQ4N32eyL1jxlmMmQRH3zQRhkmiUnpNrdDnOkacPu9/rnfZv0rr3P9
ncH0RlZdtpLUyYNuAlAZeaZhANZcZGZoEDy5h06RLm1hWQwi9Y34ZbHJZDBNjB5sUxKb70O9xGiZ
MDvNyDxkkuoscpxzmuKnhEGgfdmBw3jPi7Am7TRryrh3SnXLU0VDf9RI75ZgZi2DND5oC7asSeNu
qkAOQ+V5MBZf9sNNX+41UALLSezhLUAOrwa+yMiul8cRgZnfmxgAh8orWwjxYM7ZhxevT9ZUBf/6
RMpdlB8X6kuWrZA01U5UlmHEIXh5rFnB4pCVYiZASjgPxKPOcAs/Dee3ckWv4YFB7sOMmXcL96VL
16OWmLjbvicxWjZoTLcxqOM4vUg3TqSvximyx5D4KCWqcBNdTPB4wEcIUtYuLzJlotRlHOcOgopR
utOwWM3G5mkM7CPWQGrk9I/qk2Z/wVrKUMS79bQCzZBeyuk8555MGj8FTdMXKUwOCQbIAGZJucJn
1rj0k/0JZcigobvKY+LaFRGktexUJJKrFnm2MgF/1IcK0mn+NvYrgCSZs17H1WG936s/1/Mh06e9
btBDSqWxi5X3v7kAaVOiAOVuUzhPy9dXaUwvsEQJ9HrF1j09tklDFPbNa8zLA82CkBchSLw+wQ9c
YyR9ss8nj2Ki+0QZZl65mbJDaECdDh2sp0aU12ej3Ujo6DP4ZJwgjATW3MoqeaRKtsayerRx34gM
E9vG/WIWNPw3QXWm0ImZjWus5ZD7ujZyzUxe+9HqtGoYlmbAl/zTHLrNvXj6PKN9UzmEH2F55uyN
ywNMSmWdipVVqjKIkdQD5xUVGYyjjJ0P+915RU+xmVkf4yuOh3pY1cSqX/HIwOjBb08WM+SBEQRz
KEaiAsgQRyALFRmNaU4gnLzsjaQGgw0mNc/gjoZ1WJGWbDNIT2fATwyqe033WcmRyoaoaxd5g2a3
ta5/YggeNf03YY+HIsfAl1MX5BxH1MJtYpM7YgLW+TVeNf8y9pWNCSPLS2oAeeNsq/rwy17HYBao
dVLzFDQPTaLG0H9lzmWOI3gqvdeC/O+kQfa3UW7Y57cS2MlGWXbI/KrkySvEvAFHlglK8Bxmg+8I
tzhMXgxWNN6aZ9gkebb1pNr4rMnYUB84HaqTKtIKEeVZrir7Siap2Yf9v1bSCz8mtIV2p+zRkFt0
CmaHjmXesGmWiBlTOiK6tW7ZKYeUzb4vDs1p45jn9mA+KMrSRSEYqVXj3nUbGbS27VldKNbms2TA
Ke1e5063y8f5G52+7A1A3xB+OKGUPp14Uz8IYIFXAQuvf6notHdjbALxgT/yN0L6SgsiKxUyLPxw
P887F3fmT/zGx3Zpprw0J1Lovs4reutb9LwZSiEUwhsTqVBmOnj+ot+GxL+jlTgj+d9MaTMJQSDl
eym/ZKfNlxMFCN0jH3VfNJQy4+jvGSZyzjYMfGXlLaDhRA49xHRKcOXNr/vM/hfIEERqCnirKP0g
YWwk1grVZRG2Ise0rkRfFu9TZbF15uiDZMc25Kx9pB02/eWVhvfPFAhXMCeX4UTt3Gi0VYkc7kwe
4jqn3Bblvb1d22tddVG7hV70BrG7mTTSGFonaFFLf1IvnaPBUEhT5fhw6mmBiss1bkTxwooedC4z
sQMboNKwNjIyV2PBY9NFjk/zjz2HQHTqvTHsFjI+sMxUVlMcoumV8mMSYGfCwEgN/j/T5gQEmeZh
A7p9V07bq+kmlznDHFBCTrczT4Wyf+CYlf8lNnHj0zT2QVg+411kOn5A3LFzHpe5DxLKrjMbIsLM
2PxnzNk1MMgKrKMT659ThH1gScyg9V+nTLt3vYTPJ2c1HysM+ICtPNDuLyMdOcU2l3XoveICspp8
jZfEPz4gh3YyS6VqBgfKOoaq1k9CtttTOOAKAFqndOXmmCuLON3uaD6Uyv2dVS1yIvIS5QYutGGB
rzlkSh2M4LpWvi/mB4ZgllyyKgAhkbHkRfBBIEW+tm5s5fsji8c38hJXGTAdn5YuGE28rS4lQg4N
JRq9BFoUvQ3Z10zc7r7aJfJwsIboqRLpn9cWDj5AVgMwIrjjC1Wf+vQWji6uLgrsNTkzcSAvVvXM
x9vsjTeJvRK5C4Mz26xjDNDGDIBXlKNcb3BgdQh9erhpwr2ykxncP7ZA70ckccG68gSXrms4rdhL
bknZKKH7/vkzxXdd6nXqsqcocZypJygWbPm9Z/ZrnvZtIxfqJLYB7Li0OMf/FCcxJQqy806SFBGY
/LLDaAuh1u03dbbgomLa7ZczP2Le4DtwIHRatF9rRN3WmQ0hXgvHm3x3HmOjIEEOWebmjXCuer7A
Rv4a9ixdmBtBQpkmh8TJMyW6xxkG94H4EyXQgmryUf631djCy+Y3U621id8x4PrhVM0jkEjvMJ3c
zd28lEfjWcVzeNhlnxkVxKePB98bsRfdgxshfgya0Zc7/8BqAf0y8iJU++xkIbznf4IfWwxlv2q6
XRgr0XetiTzCwP9eKICKBNIUI08grHrr8dd6tSNvOx0Ab+yccl3WisRug04akralvAHDw7Fxb4Ek
d6HTOhCng++x+kocqSXzunkDHl7EWPPpp27QwL5IqDwZtUAKEQW26pyJ9s1ZSFMihjOg7AUea96w
SMVeEv3CWKYIVTAQVxb5XrhiZLHFuzstmthP+zdlHfxyzvvLYnBySbZ3BysNx7QcfR4Dl20j/9GA
Em8ie/cXn/1QC4V5ap3+qiszAsbQO+lrPQcY/8WdQ5//dQtOr7KFhzPcCBktPqhPQM3u/kCOQO9L
fIOfwtzG6Zi0HO2iXD6XyGqmjsLt/GEU8RGvArpfAJpWKdzasxkg0kiw3nXRFb0EYJQZpXJ5Mugr
yFOWxipVVEn1gnbBy9bb4xamoHxqhx5h53ory2o5dS0eBwCZ6M3KCXAP3Nenarxhh85Z2+PX/Xos
lX6oF9ORuiVILOUmIl33nCDg65qHMWZ6ah6Gm3y9s2gTaDoIbbWyzFxHXXMMjipQ0GVUQ+oC7TVu
i+VMMtWVKOO932vDql2X1KjaJFcJETc0yZXD/Ny/OBY7bMpefZWlM1v4/8rCfZPsPuPNtOvjQz2D
lh4fydkb8SSQNbOmRsV97t01zjSH1w5p+5KV+xiHFY2x0hScHqz1WKkHyyjYMQHxlGjN+J/Lu4He
mv7H39cqVtHl7thnTji4HpuacR5aX/m4eZ0RocUK8UyRyHDIjQ8olvazcZszpYVhoxMMEBjdlgbp
fUM4+2j2fhGgzcUca0z3bS+S3VgEzLElwt3GbO9/HEg4O6iKMxni1MHbPbHw9JWmCWyg1RdnW+r2
7DqZs2hCH36wdR6DEyDoOKNpLzEEMKfpHujynFrvQLMVnp1TtNg9gJYrXW7D3WZAJpzWgCFKzrzX
36+5Zx8y5AeGH34o6WbOTqtDO6pJvzK3M/Uwf1VtEEZpC8jt/LOKSebnfOK3yxRMqjFtVUXKTSFE
dUU/+k45LpZ28BI6q7NWY0vlaPV2V8kcsNnA5fgedxNY/xjvwH9JFT//qfhTb7FxtnsQfd0pHgr6
PtD11GxYJS6UONfpHTzWTO0xiC2qwGFWfx+HHVq112n39sJzAWEdQgySpguNqZJhf8101D2pJCEq
qvFUVgE8kitIjEClQ6E9COophAsmug5OL2nYVO+KLH6QTAY0fSXFa3CM1Cl5fBZrkwyDCIE0Yv+z
+cX9ZjVJ37dJvgn8levLnXa/Y5blpGwfpKHZKmqpq43mX8/wPHgeRAQbdvyEJJX4JcFjjcNT4hwn
gjl7WM4p+TFf03W1fL0+e8DQtAQqmAkU22GcCPpc5UMu3s4WLBE9nZyhwUcdvDkSOPIL9U6YrQqh
/1k/I/F2GhG2x/OhBtw2SCPFBAyP09wGFxfawZrfNhgskKHWHFEtTQTaXuLsLn1b/qTtQYH5Zwbw
LsdqP/b26xny4q5DSigT+c1MwIJKIkH2PkvCdPBlPdf2ByYsyh+QQ3dFv2l88qPx+246jiOQJxlI
ajBrn/F8cXAGMjdSgaC/8zAPpmNqdF6rx5fO+gOTGsbCMB+mhLsi2ctACxQt00JWGAOxL37/5bP5
ifKtfvZKxR/4d+AjFv45CgVtv/x6fzl/fb76vm4O1we9DVVe711/CnO3NGOLKb6+OhRKMMdHm94N
kh6bIRoghDx9ID5atmfW+xSVr7Q5L7hbSmOYrhLVBQkW4Y6/PBia2zELmCa4imOYTcKu0qjTfEOP
fbGF4loLznoathJFOQH8gaIirJNTkZf7exm17UeWLgXtFWCoySh6JAt/JJLQZr3TS+H+U94aufyk
HFGvg3wos+SU5lOIGYCSw6jJZ90GDLl+nN7nOvJAMgjprh8LYNKGpBPEWtEgdtTH7JFNnD9eiRuU
9RGiCeNfKk4vXdgUq4lC23FYVhzyhc6ouZ2YfuBSD5oigb2Q8Av3s4sxNxkexUFlE7Au3/ahMPKf
amlt+gzeGUP2S/894qke012Jg9esvFIVbxnNtOl74TM9m0+T+qictHmRiddIDg7wu1JZr851reYU
/q8LUIQd9Et44cTtUn+WJoFaD4vYePbIMw0HF09wywYg+38K5IhDosdkk5M+U1jxKQ06ISgDXGDU
/sEdE2T+A9Ay4md8B0IQ9I5HVT7f7KmIWFH6wEEuiLsaqK8eXvWsAH3KCStzrYLkRFSY1hyME3ZP
dt11OuZc/peU1nB4RKw7iHWirMmhd8IOqRWJuUKHG0vvJIrA7Q/uzGu6Z1osD9ar6eVR6KOZCy8M
yi8izsz4WAeR/teYx3WGTtRsQDOS3SIQpfPapJt3AD0AWwVCJRwbI5/FTa2a1VIDlVBMhN6S6mR+
icTyvKSvxmruA37H4kcGzLJwsSr0M01tlVbTaSzB9hYddRADfiKsjueZLkKF+xrp7gaB6Jfg7W8A
Of/3bibnfFRtp95EM6F4zPvATmaDU3NvR1GDoW2fOVZDniCsSegAhjTUwO7mhO5H81yupyNxcB1I
nglZQhjL75qGjYVL1K6rtcSpDzRCVl52zgdiEkf1R+uDk544vTkknecmbc8r0YPWGAG/qgGNm+H8
FfKTvcVKnAgMVGBeKb0hbkvGlqHYmzKCrmhq7L4fl45fWOE+8ShT2eo4gaQy903A94vXnETffUXT
D1l+OTgeFNrPYRlIjU2SPYOr6EJ5jCzur5VuvXoVgOrT/vxOaqSkLjrtH7z64csHXdgw2MOF2bV6
tok2OUN1hpLPBmLntHj+oZ5bCvSGv20kxQpKykGqL/fjWUDXPSo3YuUw1df074SB26vskYbkDhfe
QmFMsfKNJ/eBusgaWyLlYnTLw8T787zzcgCisfaRHzIhCvA3Ccj3oTjYB1gQFE9Mf+AtFfT3kRti
ozvnU6p2DeHxEorZX78E5ufisbSkIQkDRAC/sksta9TCig0Y4CtXV6gZdkm0yb0XUylOqTDKTOT0
3ZXYTvz6ThDYB9XTPFKy/HAje+vxVbOilOI6D9h+6S2YcxmtxPqVbwQm/HMWfjZOG7ggcl4aA/Xa
S3kUAMHy5y3pF6bT4UpxRnmWJlStjiG0eQKz0+gm/bv+uCdhNDxLBQ+Ket7Vm4nIwoGVdVbb9usN
n/Rj7jPMS6AEoh755TjaC1sxQlgpHI8kVP0ifugGd0O+ZVfr/IwN4EgQYzEv+Le5ge+SyJaOMhaE
7D2AH1bcTs4lgLNLGXbG+SuJsm4giKad6Kd6OMG0IbHs9ZYmJv53bQNFMCyGaGOR3umEWI2NBe18
IskihVREJ5jqtpTQjtEUw0UbL/v/ULEKflLjH9iKapvL+slUjcstCq4jikjOAjEJAktrndMrKFnw
3nTBP7azdHZRl+iNX9/rz8RYmVNdpkweREbcf0bDdpM7I9woMFfkFAKmWOrYjSSO8BIs3YGctsH0
AgAWm9YAffKtoewBCLlRPVI4IG0gAfnNe74v/POJjU4aZ6KeEn/ZFRSOkRjHUzAogS7nD9aLuzaL
vMYn0e+wym/BiZX6GXHQYa2Rseg99L3NplDWvndSn84tMgRF7r5Vwmbn9gAVGwJW01JaFiVJ4PrA
axGuvkTvfOviZnk9JmKN3YegIwXh3FqFOGk0xdlYJLLq+oMRTQEwfjAclq8Wt2gBTr39URJSQBNM
Tyijurz/qswkWgd9hLMwOoOj4shcCoXSM7Nmp5m+o6mLk8eLFT/8Xuobrfjh+pHBJdy7xhOJ/mxs
ovqYfyABG8NFTg1VEc447QoW17w2vNQW6qbQYy05oX1WCJ8DU3DCFYfJpQyKSQime/FOCcOpvjL3
whPTWP4ktAvfv4MqjPppMEM2/LG9IYTLYMpNNtPJkLPdNEBN++i8K/OEazkqWlTxWPiZmYYmIOvu
iQF45RD7Iw2OuzGOlAx9X+Lw+sDXGWW6cptussd+P82+4RjpWu13CniUmIB7+2pNTON0NVZtUDX1
j5c419YJTNmyQeSR5InXN3vcEic2h4JVhnEFyvNBloZC61/Ls/snRISCdsGNGnrVZ8qmrcDqlGO/
N4VrVHLhbnCDSeWxHSvIaD37bdxePN7Eowwmp/Vb4ppNLpAcb0z1MriYHStISHBCqQEh3kBBduWQ
z4tU5jYeq5oSIrNN10Jpw+BU2h9mWmAd5uryI4X6n0oZcsudI0ZgOSitlUn6Svw7YZ6SeflYd1+2
0gYdxXVY8zkRTele5F5OLIvAmG5asG3mTB3lOh0JHL71l4jzJMNhUPkT+O7sKrnsrvmGfrWlhrZ1
hPMAMkO0fnF+DweRKK5ElFpYzFIp69EN69rN+UwfLeZebBHsWMBGzVy7PnoW63VokdcqnxbxVxTd
jkzpqg04/Tzh40wiSdAPo5nGITCsChD7/+bShKRfeO04AfZe9xpC/OPuLmEf170S4oZHUJ4d2qs0
wKFefozVVX4lCTLjWq3zZM8ZDeOeorA537wcDaqhv2pATejCt1rY23DakicNGZJmYpe21uE3j755
9nfawmlVsr9PaOOjl5Yeutm0NKLoF/iUqWhEVjJD7KPt+sojzZFbkFEhbuxTsVVIDAONCjI93X1F
gMvVxPezlubbX+OXf/zVscbBKWRH91rzkpA6dGwcGwzgwX8I8MFxwUHx/fVtSNKFFFGxbClhZZyK
74WDT6PzcuyZGkJI0FZ1isdkFtHniEugEUBk4VwMON9jo3fGAZgiRSM8gyjFgI86HoZ2k0ebTajr
qOKp22TJBGIA/zzALofH9bvsyGneciI9VN2J2kB3+yDWH3U33JXN+cbhG1kaC5R6iLjcg9JiDdfg
kBXjw9btO86BOT1CFD+BulFca9BAh5u9nmVF/Hw6pTAww5cDOZ+HXAXXXghcQfuPnJGHAE2Uy7Px
44CPpw7n0jNxmTz8IA4sdRTgQ2O3aXxM7U+E9rUKh4dKO2/JIvF43Ot3y3o40DsdBcGv4GM6TjjD
LiXo68cYh/4J+RpGkUDPsKypbOETheIAddYqkwUWBl4DVxWo0H7XSyp4gvved/j8oW65PQ9MDABz
waCk+OBtnsuDXZcw9LrwgwlkO6GdVcRFIC2KpyLbCWDTQUw57/cG2VvYv8KZpf7llMawRRJExifg
X+ZFvvf9iMqQ1n6TAdIZupyqZSecaIRWs0VLHybStB2Udx7rL38jhDFwf9I8brgJeX/ZfrvE17UL
w4O+3LgFbbd0hSOea8dJ/BtP6zwF3Axot+m1PDgAxUUDbvZG3HbaTDcYbl5/NhKUrhF7yv1NDZln
3W4YhMUGjA5WXcG7nTwDRuaQch3jZR9uLFlyKB54vS5UheiwuYIdq7Udd0Qbr4LJDDDQ6Gj4nggu
L+9lJbKoBr62AAaiwsCCD6/ujmcJq7UG3VJpVf+aNIs5t3xNVOy0mQ8ihEzIsP1v5zEceam0lSBy
IKFkqGn52YYlWcH7NmPtwwG/zZLs5WWf1RcdsZ2N3ovQMZAlAbZmGlBhqSy3jE4Er0cbiEcVX8e5
SsQEq6bREenMhXeMe7o0VUlYFe3OnIf9DlXOFUam1vv5wiQqGRGTo07nB9JWm5Nd1xuiLigzw16L
o4C5dxe4Bk6F+uoqO7Zv7+ke0penX4lxYzJlZEvWAiE3BnXpRXuuOdexxq5P3kV8/fHRaCkML53H
K+dWDnljVMhDWEDTjWyfT9t/cxAinGgVUguaVRbN39fn1DyWWClef8F8xxI8mcbVw0QGRxbqgqjv
T3sdTGHsqhxKoqDGI2P7cyNdnZz951xqWgV+89zazbAJuJjXEnAwlUyEAMmXP7Cr3H6I22cXEX/Q
Atc3SBQzfYsFYMhM7ayXiwCD9W6cyIx6w3OHesPMjUHBO7E8I9tTVFBX1rEpWogQuh08ZBW1JdkU
OWeLGKx9A8/T4aa7IRIBeMUXuhU6ADfpz3xJXR6cDFn2wMQWJJAwRm6pZOjZAnBNsHSZrJxoVTva
3Dx6n1nXy1q//7YHAdmjleL3nQg4CkJrR+Lo+IAuzNxkKjb3bEcN5eDoxlBE9oLcZvx9vMzELZDI
DDMCoMvA0NBuOc04K6iRui6uTExmQ6CHy7CZOSBnmAalj7la1kec3MDCqIDF7gA2+/6z72dF0ysi
qTDfB3U5yBgPZJyLwHyRvMKRMwl+xLqfajvKUjaNHuYWKCTwnYMo9Ua4cmicLrlyWUH3S6D1aN+D
vv/jO7zWM0oRvW24zcF+dtt75bUl6YFi9Tceewif48aVuZNavqRR2kYsm3iyw4cMwwqF2LU53FKo
rMjNN1zRoo8g82DuZJF+EDU76d3rDomMgMxVRXTKI/Y7bEcmMowwDuE1Y4RIDCLMyxZr58//2rQr
CzvB+PWuMsKD6YSMS5trOiwbdPn8CvpePTKt2nSHO3/WSnNR5cmEhT4Qg9vh3FJKytrz+gyM6qpM
wHNEbxHHe2rfcYw5lNvJwYfE5nI/omkOCQtczwDXP6sDN7p0Lzjh4DOi9k1JwdG3z2cL+PC4K0+2
0Rhnaj5AGmSAPwTx38Scb4Dgo4dlOxVGH3wL1uE11afwQvLwFsKisw0gRMCpjpDMPyYnNVweO2we
454xAF3cLqmjPwmRueHHykKRpxcRDW7UBMXdT5qDY1YCh9HSfk/QD6Eya6hLbZ1C3U/SXHnb5RBn
2wjZYAR46sv0eObvEt7JlaHusK30nJSgp4CBI8DKUDaNmN2kA/l1qex0skrzO18wJkZZdWmcBjb4
s9KGWA8d/bMDKPdRDMYg7MF1rJBElEWf+uNQP2B5AaKJZwZgvAUkVLcjylhR3n0Q3LlqV/xzn+XN
wKrpgptrluoZiq2faF+OkjylgZnbsZIvpZok1gubBcLTZRcd1C62qo40BH1dOBL+V1Qw4B7U8Aip
g4S/VozUNoLFnWPD85bV9HPrB+j9pCdVhsVikIVEUDExL5FeODDkaDqXictw5dydCSX+cHVJpGGg
27b8w5nvSNpY35fk3WaaR5fmR4pww/LqOSryKHYAodM7X2QOszUxvF9O8y3d920bZJiwNrnZNtyG
Yu8M/87fok+pIdLPbCVXI+aIUtQDuKlXKhGGxVDOJqRohffYdlcxukAqkWVPKnHr1GN8NqswWeXN
w0Y2xTxQdDBLPIHG+6uQBXRKnSGcpSCXGXAX26a/cWR8YuarjtTPfFO4RK/iKEOFLwLHYdiPRptF
MEGi7/JT+Op+TNN8TRoxhFflfm42Acrz2wnzDD1PUax1azO49wX19caaN9f9ajzBuwElr726l6W8
2Vy/2NRhXQ8frNgj65GJ/wuhfv7N9+zXO2NlgnOFjQkAaF+1oSweRvU0aFVCeVvH2A9OkvdFFvMK
B4hMzxAlaB71ceJoXL0AU69E4rV+vX7ArXG2i5joR6wb3k5A0Fzt3tNidn7UMoQhUzLWqnPH2s59
P0F/Pft54hWakOmhZ0DnkkDVWdg5P1pFzUx+CsjQTsoBGROiqgq17Die2u5PTfonlRm20vd3/lr1
1SK0QV/pNVnR0LmFMezlJNTyel/Ke9KVcF5r2THaN759Uw8E00juFQV6pgsvs28ZcfCOvRv/mVqh
vQP1x2qL7pkccYLYwRSajOdbpGsgUPynz3MtV+q6zrywoBCCUUmwYWyyJAs3r7zTPjt/b86mYMYq
ayHL4XC+E7NMqQOs+ezl2X/GQsjBn/uBZNP+30+a947PCkfixmMuKZgVSzana7D0zCFMBmx/S+gx
SgWMnQWwqcba21zGNiKUxQflt3/FbjddU8aJOsEnu7IXAuMboT+onY1lufXLuG6fBV90ozS71Ozt
QvXydk2RK4YL9HW1CxjXdkAL9AtNdhqrtRSTW74viFjQYAKvZMv2a5VEWxr+HRzMc3GD6lqs9DJP
U0lVx5ok5FEzVUKKQwdGcx8ABg7y3tbTfvxDZHTsYlIzJkk6f7M0x/P7kt0TBQkMrl2oC5Htvfsf
RbiJGPtptSS3wqb7WPkDJgMLl8xdK2DfZ2n+lpKpmv0HAw7slaZPVms5CLd5UIDQlBxtFjxrOHOG
drzN3IkK68TplOBXg95HEcahW7Jo8eaOwhVuh8tN91cXa07GEH+0bsSG+7SfUqh113ZmE4JS3KOB
ih9DmmQtBEsJhQ0M2JtpS1kfvRgmifRyF11ya1P3RwhusvdGapLSYeaDxaq6U8+rnevHd+i2dzH2
7CMLFwxtcRYvl325P+ER9YyONl/qnIi+OHvvZUodHU/hg7ZntqaEDoJglYrpArnR9Obm1+zspkuO
+zmg6nidYduq1yMgKvhsjjWq2S0GtswzvfXCl4eSNKa4SeZZVMsBpb233EugropqX/B5xVjjQvXU
FhPfauRvjHIVUXP/rdHUSVIMNyMwTHu7GFgRGUTif193i3Sm6MqGIQTgp3m1IYXf1PNyY7NLzsLr
CezVLnppCAwZ7KPQz0uWIQs/0LfeKZUfRo+YY+FVNdp+i3JwGG7bc1ejOYKgkCuBj/1KB/Sdifcs
wds39ISvS43eJAx7VketB8sf/yirS5vREgJkQCLzA3x7G+jU1W8n5JOmuyx0GviywXdRB7Fl1wj5
95EYKhk5fixKWxtnOQiuTMCG9HnB3YknkWvsg2WcDHonqgZLfNb9XSFlDMngCsuTBoxqkLYIQHOA
CN29UJlHtJkqtYIZdnKaEYPGgMbiL1WhmW24gKU4Guf14r9YTf98u//VC6Lxz9GPVGwXBkmEcz/E
tc+F9qbiysGjJ8en8ez6VxFRjw26Pm+AaWKAufpC8RilPPwAHwKebLiORn0jMt6gkOf0mcaA+8LN
XXmiyIS35KGHGKOJbWUPO9csQQUrqY9b9aXFh8pfrBEAYuvHbuz2ujgNQqJZ5qooi8StZtghxuvh
ct1uvB2Hu5p6/p+0pJrUAtY8f5XHz2klMxVnD03blH3oWIITFxM/t/8mS7yk5wrKHoXvadRmbM0G
BANhnchIIYzayd53LhFk4uyU7Mm8S/054cp+7Bo1LyB8diu4VGVhDzAX86Jl6YHFP2UdnzkTe2Qq
U/OwtVEdkeTFjpng+T32iHVPvksd9ZO8Ruq2A6t0Ba8E8VeT7umGNEXlQt7WK3nhbTdQ1xeDfQd7
S4s8rMOIYn8Hx1xXFNTU2T4kHWvq5TdCHQwcWgWDjkmIUoaJa0SMzQgPemVaHxao+oJvBqsSIag+
jK0omwTWvE4VpGA9LEUU+YbhDNGdU8ZZjr6Qa2DBCgmRW4heG9IWBJJotfj3rwnGO/2rvo+5wcoc
2QXZCvx85Rh/xdDpyANm49A/NHoYfCowGfYEHVeBI5oALeSiZcPHXIEKxQls1QEg9Xpef9oKnZLd
IFAv/HaHqgeaxO4P+KD6m6LazBmAyElIvOFpyuDjB4CbxffIc5vW/B+ewW0Jc3WiNaB+5dlLezzq
VA/X+o8Bq3KPBr86erT4BbteP1Wg9M3Az06GKt532m0QWoXDNCN5T3pa4UbeG2Gv5dCvNsIy+Af4
EM8u911qqW2ZCAyH7C8slOX7XTczINeufIWP9uFK57Kk9LB+Yw9hBwHHbUMHEugXljvWgoV353cl
xoQgEtwRsZ/EcqA+wSWVCXe9i1M8w9nLEj4Wpr+KyIFSyLH88Q0ayNC91KogpOgUHb67YmZa6zTx
NOf8bS53mrHko/SfcfL4xn1i+PATSA486Nq6SlCebCyeMOVOi2Owur+e2DEYkiSG1rA2Cdrg/O7T
MEhvOTlooAtgOqN/2NMVAzARm/Lwz0nCkho6C4yIFN3SBsHogQP9A9qk5/r7a4PVQNC1u4CLUDxk
e9xTpYVWk4+W8pmw6mzf8W0Ep2PYcvVGHbM2fNMKD5Hfu3D4Wu0N/1h+oY4ihEuKexbiVE6wQlSr
LEvQlnERrMN7to2F6/mAjaUqNz7HISdpP0IJx4509Rq4W3S41BKHL0J274Guqb5PJozbRmojJSDb
0DLNUmV9Jq5pF9QPIpHlAzNw4jCXGD3gd3OrsvTzt/qiq9lUf+JZNGK4hYnVXsbkmv2y2rOT24PF
vRtseEcK6X5GA3tTpSfBcQeSw2JJiJfnNO6yh/q0dLqU5h2fTU9Pz3+IbZsD6uxROLGeUYqhW03/
DOHMWJgYmCmflNOQui9KDX/OxoPESkUPF7oohLNnIK46KlV+4QAaGXdk7Phj/DzAjBD2WSdJiXT8
4sXqXinwqGqyA/UxiVVTbbkUuvkjeIOHBavalrL7Q/JUfMRu2fMUna8kt1hiQqhfTP1ewDva4mA8
jirMn4iJngplFxYoFBPBgicm74U8rA8TFG0QMnVEf3sr88fxl+NEcoIi23t9a5dxvcTQJYAohyX8
iP9+w3N4iiac6B8JSquOMa4wrZJPznUttnr0DD8M0FTSLD33ccHAWQrT71Jnvo7SlloLMICDW7YR
6q+ge/2CynUcsSFVKkpmCJgP4MWWPnEgY69W1jXQdlMhpc94Y+A2rSZP1heDBmgJ9lpbglSz/Mr2
Cb0dW+vpzORViZSFZWnUf9TtDfh5D+8SJ3TWMwgmfzh83u26s7U3VaOWGfrgYsMbLZtUXklgmXEl
mhKGumrl85tUieiQN09J1u3y8AtqMmX0KW0cw5cduMH0Lo2zO3qudbIndMEVl5i5gqhZQ7NjSUZ3
TK77QufxFgFTZ+SZAWtLiWVWlSieZNDMuTumccUtDTcqMVpvQiF1LVXVQSd6mz7ZI3coOK62KflO
1p+6SgQFpkatvzOGzD0zgRB8cEgstRP+UddBUYj9OZo9YEZ+U8vGEV4C7QKyfUlDxeCwB1fWNBEf
mZH82rqdURNvHA1yX574rrzd3tel0tGZPgsdCmJzEWjj1NTwa/AMme+kkMvLjRMjRGLnJrWqjmLy
nsHMGp66ULobkQ4tbHb7Vdtwsvt3y+qnv4XZF4mDha3AsAKYQAxMBp8PQt/CBjAZsp4IYFS1Gu5U
k1K3FMG4/ca7/OBsxZMHApauf20dO52pd/mHRRCglGemByObYWEq6iqjtq82cWJvtbypDE7795nm
4klNgoQcgk7jIECwQSF4GFi6rg+1YJ+ty1nH4E0g9tLEtLrvICAhFJBAKDP5FqBwdq4nt+YDQGdr
ozRRRUYLdyiDjLZpNDDIoFBa+XSFIxtEFrST9J1Js7ozk3BHwONVuxof2CCa+xgjtP35R9qZ0COm
0K+ov4rZ3v7NF67SFeL76BemUer079lfPZdXO/5S5YB6+I6NbCnRdaITlQZ6fQ1nVNrze7cWYo5Z
VZv88TDJFmFoNuCNShXCAEQ8enX1PxgtzAsYxz+a1n46y46uWGjMBTjU9VT9Lap7lOOmyzWrELj5
ft2KxvlRMK04cqGWUTI6TlR2WQMfhlOmSwHcWu3SBvtCyOD+j37UvMeK9OIuB53ucPPhaCR5UURT
mI5VYd9VNbHhS9Kfy8vNXnlNvwm0PfGz5qtz0K6tOAf645VMOszm3LbtZHJmehmHTmZuDArpEgF0
xWe1P1DjkA10ZWslQm0IQPqgx75sBaZcl3iqBHdP9qTvAezOTEzlu8pujooL2PmupzoLBnJhLOIK
URpL91gKYW7vhuoP/1hF7hyV/K5e6jsyWivVpqJwV7VJvMbvFTT9RUCfKkrvCGm9pl+GR+HYUCI/
yrPO9tPxPWVzbw+KsFDYhBRzQw0JxREp5tvMbmkrCe29h1ulmg6uBL+U0D3W/fJPHXIlyw8uv42Z
6RWgEVS0MrDTa5aMPGXjdu3koWxZRbF9bWWIrddxTNlFMCh41/xIyD9JCsOylotIlzAcjxZD6dTh
hEMvYwd6QUVtrhfuOygnubATnTZAU+gZHSLzv3mKMFjQG6KFSPNple18GFwqOEMdQdMmejMVMmVF
8W4RR7z5rDHbE6v5A7ut+YzaZlqzm/afsQH4qI57ruNA+2ik3UL5tNgd1VIh5+VNT1j5jAOg/Ovf
BjmRIHeWH1JuPDUta4I5UKv7n6ihA4QhlmtZQg2c9x54ccDMKdX9emtkIEsCsN8mX1A0odGtYfOp
h3BYiGIZgnfEixiM6xNd9GdFG1JImoZwCyetWp9aklv+Y01Wo4usQapPNJ/4aW4nfRpakiQ1KKJp
HF+2ujAGW4hkdANAuq+sDsRrV/8Ae7SYulkni0q8DtP0opHmTyAXJtSJ2PGJSFR/X8YY18kPugyd
YP3T4kejikbpoWSeJ0u7yy5yQRZ7EnmJ4Ezj2g/OiY3HyQ2DKh277TmkNOuQOWB3JeB2cC7z95RP
vXUY4F2E7rOHSth6OFXJXFm5hlS+2gsLIJSCzQtqezx2NOtbCfzLhIDJweoxeu3zoN+/Es8C6lw7
d4o3WgGgZiMLICCGPRdtpppalU7ttqjgc0/J1mqSj5FLE+m0QpoF77L2lJOMHHYtNXrvQHAie4P0
A9hf021scXSFDSRxhF3wBYaOVjEstS243qYVcshRSQJMmsmXie0dyFdhXWYM19ek/NvfTLoMwUcg
2mn2Qyy/HO2etVI/70Qj+abK3/hb5A27DhwJu8y/VSErbhWOnC4kBT+QpMMiesPupT7ROQFjx4zi
VWkZhJmCZouiIBPFUFzzLuc6UCkzrkKfpaNs00OQLTyQXPlY9DpKrzV+D/Ur26f76rGYLWB6jFzG
obvBmi+Skbyf/QlNopT/UQmaFWaN0rTR4zd04g8hYwumIe3dH34lkZuqhAOaX4Zy3UU6/rCcHITQ
j4j1QcE6/7FwxZrpcW4Y7q1/UgxXrfameYRJx4iVlhbGAg3vnhtwrmvYFAnMrFJK/tvW45xeHA/B
iwOlF43kXkUESi11py1f4RAHvauZ9CoB+t/MK+A14VeVwD6KPGcqWdjbHJspbcjJdKOKAMS8edLK
K7ab7nnJonl1/xyhX/B9Z5dkvUzHgTyh9XG2sPnqICGVENysrKuXwo7rgSkXPPMOJz0PEVmMiVXM
0GYrXkh3WDgz8lcRCpuM9dlm/0qGDjrOye0J1jKWqFQh+66bcmczHF0qQoj4jXDTeaQTs2UuSg3A
YVSh2jrnq4VGSks2gwN8b0ju+VvRWNdnVwpgUVkRjHDWFoMLuoEi8xDtobGOBYJHadkAxNKAsFzp
sR11IqhodLXkm1tSLJROWOzPiVa87JudwaMvTrn4BT+FwoDuYB2elz5npOJr1UbGwQ+6hRyggxj3
MtJqN0DtTQ+Wnoezfu0HnJj6izSwwQZm1lb7AgRNwWiLRgr6hqoPdGULbz6gj07rZK0x9GsXYf6K
3FRtqwSD9VReZEKAFNnLLXL0eQc2lww/TmMYfCIye5PVvxLnnva4FNoL8MbKD0zssDP7oQxczbDz
48FcoeFOP3OKeta+7D5Cu52OL9IdslrO/t2E3MkLyaf8mOK41aItGCWikcVmMMo95+dnaGgA8SEY
qChl8V86u9nhgCiOZeUfPjpec+3AE/FkddzzRDSqSv1MuRb7a9aUqJw87kXwTODLeEnzmxT2+Sdv
NAVAN1T0zWmgCrDm6BQTBpYpRMlUCBG94KA0X2XiaO5CGfWNgo4L4e9YHjIEEYcaprGiW0bHKJuq
RleGlkKTwb1DxbRwObHS5Lw7BfdokbPJWYjBX3A49ZVkWy3rudbuxZ0nL+/38a8FcR+fA5wEe0do
CjWf/cfdaRD8hLKObS0ZzeEBxqB44jmsIYrtbEXE6pMjcFoSXluCRb+5DlDUpPiXxZVEvxUNpHKN
BmXXDFWJsrXe98z3D6NWTyYpb7/F37eC02myppe8MjShT2kd519FPfhVRPH9qJNLyhjpRsNrRqfy
oEGR6nWz1ef/RXAnGwkYuHUVWv4bDQzqmu+LV6Lyw5BIrc24tz0TytZpiDRVsr2ck74mOW7ZIzAa
OdC22+OQnErT+rD4D7aMrvXKsJJsHB9t0Jlu1OVmufDOpuDnu0YIAk4qVOUMJwHbl/bWbXaiDmxV
Pzh10NcWCRFjYqFBpPCBu0hObM72VebWkUdCGPb6pejt3RBltGkWaeGJhJuSY0lwD25Xv4bYO8JG
KiodTTl257xU/hVAqObLwTu4BWEztdnzvs23AavNZtY3WTiU8PgBK6N/9paqjS0o6CyPaisBT8Qe
3vFnz1cFKq4D0c8CjbrNvdRniitxIHZvU2Bt/2yU2Dqx1j39Thst2ATY4VLj/xYZJ5zItqAOWLDr
n6bqqWKebCjT377B0EQV2fKAsn834Y+71fOiw2yW71FcN8qPc3LA9pieMrx8YC+8P5LiC204f40U
eQZfNccWPotq6ZKCgR6B5SRzyqwHjFGl4arBEpgapF3YOYJbb+RC8Tr0NHAFLPDT8UfN1HTr3Cas
B6yWKU+NyDCLhAc1cZLn7lIqE/Ivj4wnbmx4+rdWiyt+kMSkvOChmyAsOjYTYnb5Ofc4WTiLYW1q
/vfPs0AH/qy3AgE58HHHkSmt8XzJI52xNCWGEfDLVh3Iqdwtu+ZbpE1QaaRLfr5DlcxO+wpKroWv
gdl4uWQPAuQhrUvGCjhU4jjkGRnAlPFMVLQPo6QnesTRtNqzGQgZsZtt/70pzUoluVKY7QDrcjNF
nlHjmSK2dpvLEf8zNEitHKHB8M4iHMBTof65lRzfKmP7hOg2lhDdEEuaCwH3ssGTfD0fTnYdZ+tq
DtLY+ibqRDsWGkYScKpMoMGTGNtamPrpQV2nce94Id3wABMpPr8ZoQzm5SzBcSVZwHtpkWdxF6cM
pLrpLmeap5m41bbg0pwVG7w3NulPaPOs7AW6lKYwbAry8exAjTsO/lDQPaJvWZMlw7hD6BJ/8n+G
a63Uv/QpUEFwYojJnIoz1sGZjY3lu8jyVHVcX0tu2R4yn/amH9KnQoROXOPLyIYaQZs0gwPpnzCA
XhJrPORqJS2X3gLiEo/zIhudwJlLjNusVCaERTeKaDkYX/gDS0r8RiW2Ve9AZdfO0zDZCDh4GBXn
oI4XgOpI+efjkgqmPUSUkV2g0PQS6NSObRUIzCjHeBMSqHknXI9drxmNoldW8qd73C1yXs3OWOD9
23LPotocaoxNwiymOPvrmXbAzWNNo0mTfybNOZUyX64/MG8LJgZ6ndyoebVHPzvuh/6M8kjjfdg9
ju70W1zBd9V8vpxfj2G0BmBbogZITmRWmZs4rt2qHcWCqFoKQQcuPtYowExmG+WO1VUdRW2q4sOE
P1dkuUXwJFgZRuKjEybrXxBCPrGwqv3ghA4Cj5Qtzk+UhIxFjUKZ+UV1m9z/n//iVJsubnuA90Dj
t/SfhiscmKwgjHIjaVFd1/gduKzPlIVFFXhNnFNcM+r+Bh5XAqxb7tVOfQ04bj2iP4x2LSUrGLdl
xgGANciiJdarp7gFA1TgsigzdKLxkswjEf7V7x16LB86bj4EMhhsowLC31SLt5CNOtPdA4GCBKF+
x+j9B/PNDAsut7iL6ydW/yMlXmrqSRoGE579t2jcWUUaTRGoagmIvOLdI+FsqTV5hAtkUOHoZVS+
R+/ZEfmsBOYUZxfcNi18AVJYEOxzisanlAbEYBvhEJpW5E9R3wgiEd7h5VhNE/HC5r+QJPev/qRW
usQoyK5cF+hFYLPZ/BFS+PRrVhZIw5d/SL8dAO4Y4me/BhQ4IwylPvvQdGtrYs7X6Wp6K8fEF3Q/
PSkOsKNVOOBj+fmm9CqfxE0YZv7wxcnl0nNkc4/sg2ZgnOf+DQn7vypiPEaIcbeTn450Fe5ZUYBN
WXrp/htbtMkMeNqTjF2LLPxv1daT0ViWGadopaRdMwKTcAwpdvGAhn40WV738vg3jImkfts5wXG5
1RuL8CwE+fflU65WexxK7JmHSV3vZ5J6HRKwb8aggcyD6CeXyQ+OyX1PmkPoXfY/4Wo44gGplp56
jM4DLfnYdZlOwAUOAZ5KBYW7Rwd6wBOvZdHTmMaIbJQoTpsgmlsLZfFHySxoScEnrIIRGEQOY/Ly
XY0Bptw/YSaj8L3uISJXfyM05/xleFz236u7n0qNgqtmotm1JogHnPH9zneRbWhdvzHyZIsDiCr1
o9QQt/s3islQvpI/w+xYGN3D2RVM1qTU3kjBumZCJqkbHh/kICT2EtNEdhFkQM+vKHR5fMtCcwcK
ysYL6YB+Ah9SOagJDC4HX/siblA98IArsA0QwDhjyJbKEvos6TUfU3OvEELgOH9vKb2rMDDzTtnp
2KcfIctEm4K+BpK5KvCcsa8EnCjtMyzZct/AzUY0rkZBOf1aSvfb/6uiLfRsTcDw8vTMUGKIqwux
bX+PRXoaQaUFXZNSw6iA/mtHSMsc6wV4HFgbA1RqhqQi9a9XwU5JZ4eSGlk5I1Xtxzcyt7FgovmU
Cl5ZMsIUPH0D1Ey7vIN+lmeQigc1o1reI5VD5JnqXYz7NS5Id6Dzv7g7iN9jaB3eGiKhk7NYI3xE
w9BKe41btuwkfAU8n4zkyWIxVtHA9FIalj5sC5RJNKqoGTZBjeb0iDitjb2HZodV6UK6z+HO6X5G
iGNe2latYfkC7minqkeU+M3f8VJr9g0sUyfdI+PUxU4jARcRo4c8sxQzV9kU9DrGefxoNMZcbIzu
zFd9LkpiANSYjKTzYjXOcJ9+GFymys20NuSsqP/XoRRUm/vyyqq4oiFioOhX8o0Fvp+Tu0DnAtrG
q+TshXON1aHeKj3IkdUgBGAXY3geU5uYTLVWSUX33AzXJGzyGqlRWXflwQZZAoVsZaoaaOQekMPr
rVb77gZ9ft4E2n5KIwUkXh8Wt09rp6C7CH108Uo6pHlIu1CC+zebHF+Hs//Ae3BdZkUuMZM2lxaR
qMeoV4DLJG2u7OE5qLr1661+CbvqOM8TLHTBqNJOFG4aKbSH8b/qwUQz0mFdkqckmkYjCBU2E6im
YqygfHqN3jRYoJpzQaJSo85JrJixsOQSrr3bBFneK/bMnm/y5K4BbQjfg8x0XqzkVbY1CzlPxkTb
WJdHpCF4yuzI6z9HTGWQT6X1PLPjMTY4M+VuBH1uG4YzE9xpo1HaCPJzTWxWpJM6x9IG5pFtfdm4
8LjQisl4emCrAbOYi6IOwYI35LCQCr7ON+tGgC55Emfb6rlGxbtIEmwTvZW9AGNGFadMWBTOtx/C
XlYhwJez3tkCzjcqEgRZRjMMo+feZiJD11++0fviqeMQ1tqZAXL6aZF12H/+9cnJEIY5aXJyYTh7
TYw6w7BC7/0yAbhtD4klRXzaWxdiCwK4szmpOmYVYPNUC4QRjSG6I8GQqrPIo0VPuzk/xZ6uFwPt
693cGowntk71dgb4sw9KazDX5Bs/MnotZrXWfsdPITasx/kr4xvwU1aEf0gfDEx6KYmDB1QPWtsk
nPUxqAvAVofxpAFdnSmuQhRnhDygusoFupe3GsMWZrmQvFpMdX+zOsqjifHvTFNFdjsXgaV1PY6Z
ol+9hEWjG1j0vgyhWUXV7wnD1b1qqeCazL2yb3uWfR9mknhnGfApMMWPh87Zqt7u6F9pkHIdphle
91wFqWkXqqwhnwbFndS10r2UM2sAS7tMwFlQz8X3lEAyIFGNu6OKeqhU4N3Q825/3AOUAp2ZT7CC
xFofZcPcsSV0Uvuzl26QBMxaV0CPOuHFQ7JsnqN6Z2dDVQ+yKi+woLusQTdp+Qwq0wW6Eol1ap2m
hLRmGNx6G6zNaO/FbEficMvulKKYO9ZODHVH9uzYKGSOcOS47a/Bl4kyr0OxFCYG7Lout8aOYdvI
dgy0uoAmDcQL1ilgOeRO0GrYcNvcoqU+pPPfMHAdPMLMnwpbcNhSWt+a+k9sMZ59C416ngXn4oyY
ihP3uUghR8VHqOAoX5TNGN8gq9dA0qp518OJ9/43c4krJuLkmxLJzgR+XQSXsw+GbdLxREpY9AK2
QQw6zzcI8OcADvyTSPgjSBAzlvrK2CschE7gQrwRrGdF50H2QBweg81VRFER4i0h/PHM1i2tTiTC
mwsAbYeUQSGJkifn5Gmtn8xKITEQ2foI9FYZTQALAWNTPAEayzxN0v7cI4SBHjKDSXmM2RyKGON0
3v2yEErOHSBRiFaTYcBkVax1FxNIiXUILM7qer5UOor7qdq7jZx40i3KzxdpXkOBPyLv2D0c10cb
N27dBNC/FrOdyxNyFB/XJB9JO8eRE0AdiR7EYJQRjjoRgHNuQfZ81vFOPnL5AM55lmnuaDJ0/UXM
uiVmzjm6oIWralVID/GGUercnj1bOG5laO42WHg66RUxVqq3theapUeQOOTW8ZRfN2liEpKik9NX
+veeRyun+7gULWdo7IB/hFG5J3cbaUOea3NSvvEU7iWuIgSRbEgHdt7+mgXjpr7wbTLvVfz6Ohzh
pd/t5TZgZ8TiWbFXSGrtNDlTHW79bCLhUR3RtkDBjb5xaD8y0aEvnWzoWsKfRpX+cR15j0s5Gs/M
OFjax+sunULo2D1ClKDSz/x70nZk4rJDISyHrj9WiciNqmPSrRTyyrRBJWvWGzNfZUon5H0ACfex
1J82QLnFVAL5got+MtagjWLMOUM1WTBMMawlaX5np9qDKsX0UV4WonKdMnqKw0hphM4CHj91ZcOu
fDrfwUFcCasGWxKj+qo6M+ziHXroZPZjC8kLUUfAVe6+wfvrQ2uKgrWESC7WFjF6ur/wo+3t7cwX
QTWrJ1RXAVFbVO7OvcIAZ1dEh+as4TRWkBF6Og5ihCYFYp5qcwG8CERWhrVQZBvrJcqRkvIk8vkv
N7OSq2QBESCSD4zoyYvAVwAP7Fayy9yDaenkVUNfTEnRxrra4HeDxAWQ08MorhBdBCe5U0RnGB4o
IUA4h2XpDwE8bbWUt66jK2MX8zpL6asRrTgmCCBPk8rwUBsC+eYs/burw7KNg6NtODbRDB8GQ+e4
i43DPzQGCS0+XJkFToP/UCQhqaqZMI+B03df5ERYkIE6S3bt4pQdO3SRYn0ZCeKyUSNLyMi+iAr0
dnRW46rLidyJuEA+fpRJUcXtidzYFm5WiAw8fgqj4vizYUeoEki/R67ywzpFH6tTFPayGEHZJa+Z
LZkj/+AwfS9atxeTVDc0BJMtBpJUW63GQ3Bhjtjc23CEGQbWMbmnNfRPXPZTPrr5edUDHMXVoFv9
AdtNY2EhQIkAnhAlGK/ut8J2als+Ph+pI4lA4qKV1pDwEB0MA70hS5jzbn8SAsoeWFks/sZd5ASL
83L4H45+BLO+khvh+0z8qeYSyFfD8mAnMqqfyPXYrGmNmMFpwZ47Spb3/AiigPI0rqQF4gXN5GO9
7M7dJYbknl5iRovShU6VaWvpvJeQJBgRTlGWv493UJgkrgZp3wuBn+2QqgbGHk+eBMPFFk5cKNmS
f70lUv/1fsOYhT0TYYTw+zpAWVs3JqV7IMgPuIMb/WUwfzqKoP19suUniopGu1QJbEa7wtsGgP6V
pLoGWjBk1mYEkt1ApAAbMxPlSrTRlNskCtjwy6lQPA7PXb0WakfDZ3iRJ6tq+eCuw8nvgr+7DrOk
cssQsM5AKBqdnRf7ePdQFaOQ6pnaBWjUaUhiFBdDbLOvGcEqbjOxPlg90FVxmeb4Lut8Wp79vUpX
kNlr8ORP9dPAx8tVzwDN32gZaCFDJkpEgFqotXFETDaYgCfwNVDu2+cTV8jU80Byy0sgHRcxPlZ7
ecH+6uEBYcmsPqdFY7NbuTetiYZOqdk/wJi8ymGbLUwf/xInBYad56c2gJz8A9Kf5jEOLdDVxUKq
4g9T/xvIWgHxS6s9jJa9yhXhLrHmZsoo6A+nfcPFhqr0DRZXwgqxgcwvRdaFiG7dTgR52Plg40jy
8NQDm9AFmbBDkKcBv7SSnhpb9FhYdKqDKpckT1q0MTb3ysirBgMKAEwO7yKkkmP4IPh7xHEd4vai
lJat2z68oPZZGsXof3uvfDes58w9orSjs7oAIxNvT6a6wkJwpOsNicwdLpmta+FsOC/qLmZJ+RSo
pVjvrRiNIoz65FYO9CFXCRYhgayZ9lELIHZEjCRew8wufVRCfwUGhNOaY0O9WWT1ZE66ZxsXz8XD
5D1/9bKk+ULDXapJ+f7KhytaXM2thYcmN2QbCC3VDthau+x1dFSUrqqnMGzae5Lvtqe0RMHEeoXh
gT8mOYrsBNM06jKjH7/6G9J09f9wZVchxsctIdL3/Flk/OszpTQmWwMTP1y2Wqqft0+DT/lw9Hrz
7Tib+9LFQhpwVkZsI8x7EWIaWlzq4BUjfS80IZGogXgihlZ6Lxku68BSK4qtSBkSTRddlfuSveK0
i6Sjv4iixwn0eqW7lQbxwJoKcH8JuBQGSUodwy8CcX9Vk1Yzs7CejMBF7+cjGWb7L8xH93Mx8DsN
wpJ0r2iNjGJSgN/VoF2FW7ld19UDbwsVV2Q0kYjeAseeDX3Sunx9E0iYTUvVMHOgFgXLN0/RqqqS
qhnmKKRPsEjqZwbOgzoMLaeDMp/NaEn9QKIDYJOBmYSJuSujIREaOa2UN9gfDgtc4lnYA0t0S21y
EJuylpwG4iL/FPqknbQrfePQ6nLchwm3DQBbhWTzG9JXYZKJ5YaMXaTYt5BtNkicTlVspOj0lI0f
8fxcl4fg4UyIS3M5zJ0koIr9msdVWyax01c8F/XiAD9bWFWFiU45A8401f1pRSp8TDtANqgs1fKn
WQRmQCgrRi8xw3sfSoyvMqJzjo8baWHGRVFFYtUPPOT09imNHV5E5nplXYSz6Y8n07ECzBETHXsK
qkje7ctymDvtNYb1iDncaHBrLD3Zxxd2xxwtwSBozwAHtJvyjodzQEjn9qoRl4Ghlt6PhWdkIeY1
bGk+AKOLv+HZrAPnIKjWCerhYpAQrsr346FBTgl55aZnseNT5QVwcrirM50cjWBoW+1XG3dUXyQ6
jRJE/hNGuleBkTmv0tKop9EmtrfHY6o1EmCoChHXpttdKbmoJw6RYjSPcgppQTB8fYWyYkjZQQRc
aWgKeziwMWaogYXX/kI+ngVLJdlv6bXWlIBEsEvkW/OOWyQ66PuiC1MN21lKLmMgZKddrK27R/eE
0HKnluEUlsUmEDsOJ96Icaauf+95ItZoSXyjHxmpZqVcOhvPrUAbmoPusoarF+EjX4HZPNsrjnBK
w1rXZlF2j3mcBDFqwyh4VHD3yA5s4L8dhaKZBs0HcG8FoIVIC1PQk+Qlo85k2RBhXFOivaEqU0ma
DiLEOswFHXGNaMCcSWjsk4MvPJpITCBiZansSptsMdTqDCpc++52CgZwNHzWvXpJZNg7E6rOp5l3
y0ooKc/cbmiirYfFFjELv37HliEqWABKBGlMdyq/NfgGdJUdB1YiG0G7BTpFsXmiZSKJ3LyD3zm5
vZsnrgxDV63ZljHVNX+G9f6WTrhSCHKZ0RoUMbhIjEhfnetRcNrnV5m8FiaFUHVSb99nQdcvosUe
JQHilYkhQZODffURGw0V+xXFm5yGsDleR2hGETELtsZlKbiTGyP/GHykfbhhbngufN2IBm3kzBOs
xz1GqLvWHX1xhBjveDcR9fGaNsp3oEXn5WMoK1knuyliq/RNQRlLNrQwFxSCAB9TuIhJyj5MXfEf
N4yUgyKJLPMlYbZEXvihFjp7quMsK67bnSVWOlqrfs/gRcsS66w0b+Gs6mEIqWCVfYKAWpFISSr3
naN/gX9fZa6/XLTlxqYW56ZJJF0r3YYKziZmbA/mdxyf1YKIWL/LyJyh05rN0f2UFdCpAmlTV8+a
8iBgoVAMC7ehzBx3MqcIjSHmBOUomD7FH+w+h6LKOWrGqO7fAemV1dQgqqRy0+ysfjZG1/zhbXWi
U/P2WIB28sJTmc9N9XsbJQL8cD/5KJdoaP0z+hB0e8uOB8HOSGuNYJ5JEHDOQGJXeCdvrB2XNsLt
1vd0AiDWujSv56ZjookD1tsqal8bdGgTKNU7RaeoytfXy0fNmBaYFd0VUJ9nPk+LFipUaUTuXhEx
VtxP/8EOwrz2g8BMZj4UZB0yQPggUj2TVFCuXuBVxyABRm4s6typg9sqrzLdpuUjgwIAE/b6kED7
+96bOsXBFqLG/nG+ktWjqKNnuhk9Ua8okpSlWPaC7KLo0NGbi1mtZjYfBPEE2SXrUUH8XsffE/MQ
icJwYbwNeUS0WveSV3DA81q+ZJGtNESMRLhSbFPNWWta6P0sgxryDm9FSbBPKf6A4iEDSH0tapPB
2BXpRPWbh/5eLHBr8R3ExA4IFiiN/EJW1rZpd0w0zAxofl9T0axH0dp/1Uxg1yjt+AzavYm0L+mO
lP5OJS9gnvIddugmGg11ET7Q/9PDYz6penN6t6uqn0tkuzWmghQ6JZgJ4mXK3abYRamaN2D26GMR
7k+lwYyvygEIu+3Zydmm1GKutUqS8mEv1ky+SOiwr9aZ1MDbTZRz/ekvv3A5ugwiRlujWSWz985r
77/Miiq8kEwN/dgIcjwkcElhwCWKGV2U9yhDDo/v7vVYEgfDhxhyakYU2PQjXvT1l2TeB2htKUFU
ZWCMyqydJlmzqDlNUWEYdXomu5hwCT4PY6bctiklmeLdQnpMOyhDj+/2h+++7sMSF47fso2t9AUd
C8OHswI0htt6sFKhwKQMv9BpabAMgawL6GZJwiJFuvTBZr3xR+fWxtUgHRG2CaI848xaI5+2Amoc
Sth6jTiQt7ERdBkS1aME5VJguslW5vFUcEJzdIg2XiTK7V07U50NxFabVlRVD6gvv7mtu/Y9SkJN
72nllCasgJ70ccmcjD4LaUx8J4vG7h9XyIlKHoh/nfYodiieYYjJJ8WLcVDLRGG89dSCnIvIAZPK
nKjUWwNyV+cZ44orMH5Sn+/o8kjzlbTflLd2a39UyclNPuXjej6xRuowJNSi6TtRZyaRR6JLSWhc
H/wPijEK7kchnp6ZVrmejs4cWa39eH3XG8UxxWqauWYk+5Qnb5KhFBT/vKESLbWHFQ/5IxcTg5Oa
6pogY2UQixkRrdNSfqwrFy7vT6eCcwOTpuok1lNALvrwr5JoowvfZi4KMSqi4Osla9DQ4Vwg5llK
SIi0r0bAksOKYbJqDHJwRk05Mf4RLbYabt+vokPs9u/iTxTiQE/VWPlNkU/kMLQvycue5pBJOFsW
3a2Z9VwBD3FAJQpkugLSoFKQKdOdV6MHuZcuIjDzc5zu2ULebtCZSh7N6Z8mAkmQBtWWn4V9G5VH
dwi23F+WGj06PSSDDxSZc+2BAJQA24+W+8YFscm2UY4YfuNpBRHKjt/w8O5icGrb7vFoazWijOAq
1grYs79/f1GfOrZwCqAZlFwVIhtNj9pDqQbmhhJFFtjcHqbHTi6Lq5dwVoSFrAD7rTXP1sVBZoRg
aV4jy7Z1eMZP3YaWjZPMC67jtsJRt7C1qMYfEccU5BASxeAVA1Rsu/w0DTkkcA7WfP+8ecaWXRJJ
WxYxfA9Znf0Zsj9a3qpBXvvSxSIGr2fF2tbSpK0PQGInHbEi+XqaR4aUrhl/SJrMhyVT6PSYyrA0
f+/XZ8TMEjlzsUQPQIpGsZvjSJg9lDiXaih72Lp+TGyGP+w4wHeGHpc+gGNzGBJGcF7bUfpp7b00
INT2tbsZtSljTBEUGKXMgRL3pF4XPxUJwHO3Wg4YwWDigAu9xkr789eAkcNKhD82rwEUltkMliuZ
tivd68flaqXisafB9wmEcl02IsI+KmkhDiXAPVHcfdSI19l1fcX29vmN8LDvE4czewjGKdAuz02S
c80xlSWVS4eAMTMVBgbC5kToow/4Nx1o2Q9q6qU1dBC8U8L+rdi4zGD1zs11pcRbcXXgYOcvM8b0
DZ0EAGnFHn9/RMGso2CObXJipXYi9BjI7aYgcV0riUk4qvRvyR+AU/VPDZ4qHAC3+cMI2VPNdL3L
Zc43LvTaf9H+6FSYQ+zl/Iks3wkdDIBzMrU5ZF9GcNOrc/gKlxSMicNcXLakadCqCTuAlZRpbmDt
MK9e+2nqOyA7/HD/C8cxrLJpPTzBgqFfLRCXGlalAC89ExZQD+EHR912R11uE4+i7Yl62g9FbamJ
zQvBh7Hrc0k0PYH+jUdfUUOKOaUUBRjDW6zLYrY7qaw+qZNxP7akN3+NtBqhMOjGm/U1VY/py6Rm
E2UgqJ2yi1d3Z/lCGUQ1kgbe0PA7FtnJVnvxwOk97zsAMUxSbqey2i3UY0exapedSekDQTA6mwQV
ErRUKruwJKn6hGKNUFWm7YDtLfw8L/kKyRHWgOGZeuTiFRmi5YEY+/mjOPd3mLMp126RGpXYtbP3
HW83yLzjnfjDh2eqUBO1LoxHv41TdbSyY6P9h6HGcX+5Ue9L9AsCaLmzMeLj70G6j3IzmRTNue/V
47j/VmadB8nu23/+bm73OaGe07E8ZUQDhP7tzfXP19AeSZDsPZOAsnTtf4729uQts5lP434r4Aea
LoaLYiSMqKSz917nX2T4ULTr/ATZ+pXtQyBSdgKetLAi+Bh1T7V5Uj4sbpLvx7xQofvwpq9SsI0S
25y6GSgCpcn51sA2lKd+Za6IhEHWq5LEZy6csjozWqBAJXWG6ocb/knecUG21oUUvd7X3BzlYZWS
UZQ9VkfWlM91eKTvnJE8/4O4faD+NvIA16i9G484LXqUKVSz5J6R1Fc8Gxqw5KsRtR95sQLQJ0AM
TRNZLwTK8NjWcocp7WAM7BcCgsxsJTcrJNUKxvJYDv2oONEHeM7G3QMiIE+wz+7B7TRGWjWIoCzS
otH+yiP42TgOxgYSY/GAv0l18XoNWbsAbYWZB4JLdARtf2HtFKyWV5/SWJFV76KWz1jBI5p784Li
CTjj07LeoYdeeFh9dPlsrB6kw9xfvBjDRkyGdGtLBF+m5Fsx1bOIkujvboiXN2Dk0daFcc52giZC
60e6E5GaeKflyKRK0bKFJhEmjbfGsGIuEqGJ75ITimwJXDiCyqucq7tySC135dZjEwwO5OJXgzP8
eeY3qCSOZRLKTN3c7Oxx8oXdi4MiQlrKWNSBaRE8DJoJ3mtHMDO62SJnNmmjsVWnPpQ20iMidn2I
YTGmRYiGTfT0Kxuq9sy5XgHdpBNglbCgCS8XCdLA6bsZ7DMAhx5rF+oCba+tLkP5WJiRcYLRdUjY
rQ8/F8lfre64NHLK3iWDO74STfRy1c3Lv3BMqLWaZj878K1EJ4DfH07Pdh25VfADt966xtPPEZqs
AaxsgcoOGEEDRJziDgAf6/gfyAH4Kq1hotmVtRGCUCV0UhVEvBgMtJIU3jDmLAl1tmyypANHN2J5
94TCUjsLu5MCp5fkzAEJLCV+zVxcGgosaWtMZ8oi3rdgLje2CN+vI91w+Hrv2biOmxoy6SGmVSdl
zMwygAaUcasVxvpdBVLyL77vCLw+4nTWK5Bmyjrha68Cni/fq6OBRyXS/NKwkNIA6fKz7yjEJHBH
obCRqzEQZ9NPpx0hq9SBcokLN68W2sF7SAnSM0qOLEMtZHeYnAFn1EQwks7YeQ9iSaITYkMB/iCZ
riHfgqGbscTFxkOt/Fs0NbTkRyo4RG9CtvcHRd2dbA4AZ3jZu8A0fRlAOqiQPHxEJi90QVtP+RPm
o1QZAGnZGTcdywfnnX2spyNJgpFi1m4H7qRra0drKlK1YgED2fUPOEpVaRyY1lKFtTOlcNprFfPj
aPRK1Y2ngceCkS/1Zo1ZnMNgsZMkmzFWhF33bhbPsuz7OlUxrp2gSXQfyWiVziw+tMvWzZiwO0Vb
1lz8qC6svFi6tkJwQjF7QcYP2N0SEkHgRxKHv/Dg5hK8N49mWxkqlPhyTYnp+Fa1z/Vqobag/nDF
NWRmXtxnRxdY6qAHIYu4E76aI08Vdbnf7p8RwKBGYLv5Gg6d1Q9ZgweKior85slk9NHlYxClfHie
wlAJdTK6KbTiQmtCV5ad9MqCuprZzns0f+EpGlFh3Lbq3ejG7Lm6S8g31koDIhQixsLb1jJg33MX
4PhjsxHHsQCfPaI3xsCoJhY3MleyU3Gzjm/JZcQOuIJOhfZkxcZdR9wnEx3oNyzsErn8FDUZpTY3
p2yRLvAJ0ogkj2qUvZtxIyWol+NsKDg/7uzXh7St1bR+H2/HGxK2PhODMUurUagwQxXml2MEDwmy
Y5Iuecv0E6L2eONWFbJeQ1dpgIDpmxrIza9nSo35PilcYWK/gdFAhlbC3omN4feYR9OTcDq3Ihy4
r7jwfE1Uoq8chmwYGZJELPtCa5AHycP5C1WKUT0a74lCG1xJPi+0YD5KyPrMPjohx/uQD4LuelzH
yQTa+IwAgC5D01h8VDmA/AH/crOCsI/05W3gm5sneISBu8jGttf/07AaYQBCeoDW9zHZujK92fzr
riYk9yn8ShbD99V7LPws1dILhhs7LUl0PKvjPCRw3OqsljZaw09ICAv04dK9zGcjMrbJ8SmzCNSg
hlX/SajSUjVhCVKqKML8mL2kMTfPYcZKa6iJtgq9J/D4PDh03UodhfhiU4axSJnqwMuYpKLCbLsy
JrT0fk5l5mXpvgCdma2szzw2kZArVOclfDfgUdRGctYZNpT7XV3TUkrKpOEztJcjdYAkoov7ohDo
1FgP3667vAt0jn5W+A0Lj+Gv6FIPp4nZCHmP9RWorKsHvewPKCvyMKp6T+xuH6I4jwvr3Pw2UHPA
yW9jO8HHg3/etkHce8eyGGtbhxdOSGnRY8tWWyXyCpHQ9jil3MY0RUXbYkRTyeqTJTTdY3O69mY1
XkvRfK4C0ZPvJTL3Sr3VPWKr0H8eCIThY1Z3pAc3Ck4rLJtl+RyRuek6o3nl3/REoYRGFd1KFvOj
EAwGn3g3ToRmKQbHnfa+Eo0dySCtMCmeLgojjpbzmhpGC8L86buW/54Iba98de17es8qrP73yqUZ
hDaBrwknmnYz85nLLYu3TWW09J7I5khlAl6/rEUu0DKxhuPZQhaH7BRqUM1wFGwrUHZLze9Sdp38
HrR9WnPhdkt4dp/GqnXtMHrdQxCY9V0j4qdMEyErxkRHjXbLMR/+8xPXZLx/0UkYs01BvdmN/0T2
NbTSB4jfm14B5KQQvMu99TngpAy6be08a49NWNlADssfJkoRtT6rLQ2scklpen8FY6WxtXLWyU/F
xn6EDckCIox9xr8wkHYSHdaSHf1JaBz5ScV+ebP1z3nUF+6cTPUPZ2AYTOXM+61uucI7xYIuzl7P
+twSqUXlYnxkELFvVu9rci/+5tSnBa1w25+BVGSCr7JPPvFO+3L/divsAiExMFGGVDmoWu1CFFkt
R6A46gqVxp7wqNNHUZiYl1vrLcx1zuCoL0EFgYbHK6xlbVQZUIFus55t+ZZxqS/alPQ36CoJQTRm
CS/tq9WtaiHQOvZ3cv2Y7/iAlXJkjsVLuqghFTgjBefblbEnHJBZ+JNWeiuDHuHUfg+4PDQbVzOw
2K2T2HDLERsJlIJ4LiwaXx0Mujb/CGqkOTOTEA0VNWzmEQoluQp0cqaQiX65ra8xrT4UwbRUdjgY
BjjCv9vDdzONxiVWpNdTwWiMzvtk8wcBd9cUG5RtmTBouprxPQ1HIzdIl7JXjpzwp0DOU5q8VV2B
A5LhFkrfgxuWLQVOGYJ+2D8dhsETdWCu0b6Xob22L91KuyGDgzXY2i70O42lBP7qZnkSrEz0zOpR
xzHGqlrScdxmGqnUC4ACM4wBWl36rV4iAe8Q0MTjS7WxZnEX4pVzohcRGBS7yQVTcRDIT050+TNS
F0Jp5m7AxpSrMesaszMn6DGVmZdGspTsiieWmP46ETti3RTJZNBG+3Kyt4j5yZwYECYZr5DVAmK7
pMbbZoTbcJl+NWYNeD6Fa2TlYpkQaPZEUx2lEiEHLo1o9FskG9UwSpcfh34gnORGLyQoLbpoNmms
Ds9PCYmO4BxUFcFBGRG/v/fCOdHyJE2KxmAMlRWOeZW6qWWGXU/nIFS2pN++tx2CeFgpi7n3CfNQ
vSKvhSuWqC/KuQ5xXgPaKEAIHyBfqz5D60XRJ2dqDNh0VakVyE91cZfNUFLo8mEiwM72zpogaShp
zRo8WdvkugbmLZx89YHLb8E6RkhGilnhIalJUWMOEgSPIFbmMiCVkhYtE2bCN+CepFAYs0jW+D1c
fKjCyWn4US40tgZarf3I+BQUDeDZGm8m60aLEotrUbpYjIEQ0dDHu40ME86LbEJii1w7hCCxF+7j
12uVWvdD6pUM4PENFHYYlyo/VQCu2lZ3rLUAU3sWigB5BkI6NWf7B1xVNh9HLxKMgdoEGcDgqW0Z
Kh3wmzsK1vbMqEDnsQSSBCGIzr5rzB1KmTJwAlFPjR7p2jaEdQUDDBgc8K3fb+La34Qe41JWOfqY
ql3uLZNMWWAPPFCEKhzfIltUCDuDoxPJJZNSmYDK6mdsoXAjs3mVO4m9TUojsksCyHOQoQcmeq0A
6cZePrBx8f7WTQ6lGH1XqlNmFj7lFmPI4ioFJx4zODTSgOP6DoFUgA1ToGtuOM0xULDB4+haWIia
OyzXungfwgs+fghKJwBMFYAVAgccnjQDM8qbSN78UWdsKYry5e7Df2ritGJNqT7PJbJ7ixjpWtx/
y03c39cT+nNES1yClyVcmNT3z6ksM18Dxtwc8NL09u2mws8UzRHc+qo/9dLli3BVpptSZJYAuN7a
rX/vzwxpQ7EQ1aIgPod9T4yHbixvlvudyaIX+elFrpCsh0BYYVECy4pK/txn6ScfSEejiwP2UNZs
CQYfm+lizdy5inArkVXyqRYtjdeQniTD7cajpECyGiLRvtQxMyY9JpeL6spRrzyAMc2aq+CNuEnl
ciJpgMIbA8VhoD583vTYhOITMuqgDVRSSiQQfPdGmFfhlE8hZ1rrggMqKiTpkNZpptWDGaiwvcm7
KaEzXIS8Yly7miRGzbpoGDg4mmzJneBsyNUzNYqOJDfkx0NXOd4PsC6Cc0D7Y4jw/2QwMOnOvkUL
uLGE8u3e4oeGvbaUejiddEdJ8wYej9BnhqE9fK3DOMavosBq9D7rgE0hZprxXlKUELLxfTeDO6+9
51DzVTTpw9c+Y6j6F+sfKFGXRL4B3QAg9/lUX9d33hkYTNQlegND6nPKRv0eQDX4cp5GNvLn3NFe
+jcCGMGdiBXCp1jD1TaqrPL8iCHc0ONDF73JS2v3Ck2RsLE1nUW3ZEy5YJRq112Q0eSnqk+uWEf4
A7M6XK/2achv9oMIGY9NtmaC8CZEJRE5EKXpHLIaYeqOl9nicn9j2LWgmebjJ9j0G8NDNOpf1FJ6
MZ0AcsHdWRwtZYf8B7+yyJhOKglK7UtfPBcs9iqO49O0PfMTFDRV1UKDXqbHglrcnO2lT8mJAKqi
TW3AQihL9X2Vi+WWI+yr8zAqU+3tzCRgFLWSvkuLuFKUJtHP57upxB8Rn1Cy/CDxvGkAVuRob7RX
x1FQlwlOLieS0TlJ6kzdxw1JhsGAFhPCbLHSrFJR05/X2LkG8//YYmwQ3CzhZTzynxR62XYa7kmi
ZeaxeYg1CQLTLK7N9SlYndwcVMXHxc0FWJ2WeYTdYJWfODgNysV4ei5sWq/jccFyxATzOOa/G/VA
L8cj0NYnVT5ZnqNVaL8Q5DXqiLdhtX27/qv2m2R1wFv3w8JpcE6c+AnHEVDcnUm8zrJBSXHpk2j1
ohJICMCQYpNP+rUUXJEJhuRQ4MvDy+DMCmRyXtUxN+/lPE+V7VOtJGMp4zWmJ2X5Ji6undyewMvf
Mvbjt3AAitFHLnt/uLzcttJ+bp6RyYDeb9GUd31+9tLhyxaSFyI0hpgrDTjcii7yZ8yk/y/5MXXC
0N+iMXlHu1srfFOfjDRUJ/VnsZHlcRXlW0umdM6U6uMChZoDFndo7xT2G2YVTMIyJmjTcyyKgRYv
w8P0Kx6w0xA9CkljP899kD5yB77PoAILG4lQiWm/E9uWtHz8TeL4Dun5PegKhhFgR+gAZHErwlaN
Y9Thg13iRozge9cYt5yQfVAn12M3eJI8cWOadzh9zk3qts0kDv4nyv3gC1e+3+9Z0w4defZO0T9Z
cJReo5OtSaiUeMZ7BgH70b5QvPVo4S5kArjQ6TqeVjaY2Yp333epLigrSo5lfSq7eLD+K6czfQGq
Dqg+c8ZboWFQeL0aFztYp8SaMUo3/N1CKJT/o7lhi9NRHGEcpV5AaSJPkuiXeYRuijNoPpuq3GbQ
FubqhIx9QOp5pSqQG/vAP+XYPgxsAteiC+x3RPCGqsEy2FErrSyPyPu9EDCzJMdB6Fwt8Xx/p7tq
bbM9FMmDEk+qpeG2/nUGWTlnH9Xv+BFSCbztLvtmA7gl2USl97mDaRcbmWi5OmiJ+hPhLpX+wLHf
RatvIYdrLsf/shLibAdKsIChF71/qr2/MoDrglwqe+LVhvSZYLmC9Ih+zU1I8NOHfhmHL7W0zKYK
1Zq+3uuTeHuvCrrhK6mztfMpEhTJMbO+eQJGVuWhkeJAtKGoXvr7RYY2zrSLNAdMdiUZ/8pifdEO
OsQVikAvdydPpkPbK2HrGQuXZfpF+Y5PZf8lhZky57d17L5y0IglUgAksqayYOa2cFu0k70a5k8N
1udF1PkkStNJ8CjgA9Do908c9CI+IoX5IsO0Baz56VVqXsao1MNbhNuRW4qKfEVwZzJbXDxpzVrN
9Ec7faGlLEkpMiYy3uWYnxfZT1GhnFanIP28lYfIcNSmEt513DUqBV7bUwpBic3v65GMlIhRG7jL
cRroUpLJl8SpjnbJxHtRmUrVHT123xismLmjYoGNYpwHk4HN0s05eI5QilUC7nU17LcqLjFEcX/z
VAfVgl4ahzp6tgXEvjgzHaxLE3o0/Yrxt08A9iWS8sgAOSD3Znn56g3vgjATwD7YDrjLrP3s3Het
nSRPHC/HAXOg107WQN/IaOeUr42VOsvIZX8Jjb1Vsw/NnziH+cmK1KY3XuSZYdIHUiM01A/p07AA
WnBAx8vP5Wt3TfSp9ybECHzFiVQYO80xfg98Z/n6mQ+skhHfniKFy15yaCP67aFQVmej8572aImb
BINbsAMFsjRE0c+XnuGfK0TOP6RBNQO2RGKEFnvQk4XsvbGE64NTLqHMVdRVN07nkQ2deCgIO9M0
5YJb+SVh9w27vYHfohKkTX9xol34TIhBLXgbXwgUYOxDtHH3O/f+HMmBlmE+8b3B4sxRa3t7vXnc
ewN2fBYyVhHFsfO1F4sxfM/Pg2jEtGz+P+FsxPyQ9WqvcpI6gYwVwv8YKgNwxzoen7XHfR04Ed3O
oW1RYxoQMoO+MWlLYUozBU5S5IZ15J26M2E49dB8Mhl9znS9yQhRHhZREOXsvINJQnWonOfpd+Z/
+csq4aEHNC1A3uXMxxDX44oPSTggzHj5eXzFGzhHztlHjDp4kcM3THOjwqnIBfeMqH+2vRzP7MhR
c72zah53RdHshcQKvxsxUISbSk+aKw9aV7alR/ds4aeW66W2oC0uiGSjskPP4UDj53Vm3WyhJYMX
I0GOepckhcHl+t+7k72aCfZoYADPKzazNgndozupbc5COu8eQWJYU0WHDHEjvzgSxcdMO25uIDNz
++dnrnJeIbFJ5UwckeyUx95V0YIi+N5hoRNwJzBBUBr5djo40QZaQVnSV2uGoazgLRyfO/DIVG2H
fIWw/41h0W9X10VfSqmMSDarNiybGCnaaWx4w7qyugd3uWjW100AzQ678VYuLy92WslS6Ywsj2Dm
AlWHCtSd5Gr/tQnLkJY1IOKMRG2KwnyClK2i6dQ9HWWByb1SHBc0RSVi1fffyqAF5lpD9off9+Bb
IUEFjk9zLrSEPwRZoLv2CdM7YzNtxHw3umefMllykoAtAgu8F8ZT1N7CUsLltoYI0muWmuJsIUAC
jL7K85gDsVhmyld+74JTba26lxs2EPCaCmATbxP4AQnfeOn3lfc1ntLgXJHk7mA7Ucbt+stn4q/r
ktDwyGp27cthKNj3F4yrGHjrfoQK+36Y6kBHFdxDujvWu0DqmLEORWZtuAiOa5hznooDd2XoszPH
mWoAM4Z9S9FMqlPFf6ux5C9YgzZjiySExX6p6Z3Sjk6tL+rTdT4dSc2C9mn9JF+pV8NauZv55Woi
xzvOTvIQGOOQbX9By4Z/KYoSpHP608kiKiJIFicodCSdwd20tkxUok5rEJ9miAM1TU14TVIHQbqz
351uG16qoqxNtBy5cwmQWqzl2k1BfObL7hX3hmaG4DvE9gJaKR2r/X71R7VLjvncfoHS1kqcJ3Pc
gK2eEwghwzYKa4MzfMZsWwiQ98VhwSF3wArxFHGmQ/54ETXGE0YTgGxCpfnfK3PMiHMRkbwAkzc6
NObXGTZyJNeqVyWSsheB9hleNwFA4O0NEcz+rFNEWgkQ//NPQtRiUZRnm7KEeGOai+/yMpblGf2w
r5kbcjqY/unYRFe8Ih/+RkIyA2tmp8FVzJn2/gK7n3snzmS70HzWpQDdS/p7JJXGafRnSAfMV4k8
1Pr130V0+L33Y+xSqu5zFkYsvXmbFTao9H1IFrDaBk1eyy7CMY2MfkglcjSIMnLo1TVpgrIrT/Nr
vmGqjqhM664/cIYZCFgZDP5Pl2FJSB3okVjwYxK4wPBLl+fDLrtApyJBiDzr3vBfiRtBnU63GQRd
HqHuT6Uc4o8Ai8Jtn55TCFX+uTnWO2HI1NgiAtTJy3dw++PnE3IvZhh36VE6aCZcUYL9CHfHsvsl
Ukm+vWOeGXzaK4suOYZtLCl7/IqhkX8G7pOodoP0I8QBwk7y1Yxp5N9laARhpoivdTkApdSGdSKF
/pDTCJmL22bDat5PKdkWfez4tzWAmOtBeKP15IDXFO2ApaT5W+o1Bam+smNIZDvUXY1jr8Sal1XJ
7qsW/0FkLxGqTFGiH6QcnMz90c0kUt1Ti1FCmlMUsEAv7kJWqLuXe5Dzxr+60Hzp4GBUYAj0s89u
NUsiPnoVwyLn1VflZho0Yc/4D686FKTU3+/blPT78AT1Qj29jiga7/YP9DOC+VU6xdIWo9WzblZG
HiopQB0RH7/iBdGxi8nYIUGMKOgNpN+evEeN1uA1NIHUTzmsqyxChV7D1zND2PRODny7QDnOaS42
zurbZV3hfDtLstYSHhzdaP+WDxJtQ/ftv9Q9tQzTjxW0X5lQWA0S1c/BXBC+fpJ1Ne5zubKd4XfW
0854x6k5uOdJ9QUNcQESWQ75prS9YqFxpl54Yp7bxNBYgis9e2DR+XAISDZHm42SbF83RYhn70ms
lnMD9CWJm7uuA750+3sGgwIv/3bTW7jDzJRsgQyE7rbuJJmTf6FkE4A/BQ14qoTIZaK4Oxj/uGZ3
rdSPEbmr1leHr7m4tk28HsFOgmjTFb7UOW8bO0sigHSBY3ET5JIgqpBxxJKe0+WauConf2LBeFLY
SCthMxtBF2TgEgzd9KdT2JzEoqezBaVLy8WMQiowcOIWmrmqRHj9x/2HXOiLInxgggwcz7195OBr
lLsA3gLs9f0OLJxuOHvFq7MlsoncK0ycd7TTjdxOJdNozzEFJPudT+Gtbibss+0GCBISp1UhWnxn
rn1faD3LTeFbPm+p/txqnegnEF2Mk08dgUg3dU1hFrd+Hu6JvIV7+jBq4+qOzYdC2VLsrZh1y+u0
xH31wBIsNMVg/ThKsUTyegWFtZU2Qs1I8w+2REICeeSqTWQQIymcI3YW07pgv4dq3EMb2SzG0PMr
PwyWKAKl1z30rvxmDqeMvc8mYWgqnZLWK/XToupirQyES6IqzSKlKP8PGG0bwNOTE6SP+2DeTSRn
CfaeRFkGoqokhG6G0pyijN6apZxPF4tR2D2CfxPRP1wYbrJIPukrJyTEGyHBikrWubfrsv4jX7+E
wdT4hBOGZYQCZJIGrSiHMsdBskssDUYcxiDJHRVCcBXUTPA+YOb776NkJIohblvrph/AF+SHGXRj
/ypUZq8miR//wAof7tQOqhfS6LVlXQOOUpNe4Fw130MTbWknDkJh6co5IUzTHKSt9n2rKY4b31or
ksa2HCJ9JJg3OxD4ggrM4qGBSMAbYNyQxKyKXoLvOtT3Nhk8yuoadzwQ1tTH6+s12gaoBHEM6rx4
fqKxDCcdLbZgf5mNmDotzrNcCyGZ7q+aNtn7PoqTGED8ppChK9MH/XQS7HzJi7jbCGW3lnadP9df
4Pegi9Wfq1i2n8uYIsa3c2AP56holHb51vrhc40CKkbJjU/4sFpV9Kq2IEKXftLgvYdQUYs9942A
UfrgdNXMyUx25ZCs6VdzNG3ABAp8egQmIon9W1hoONafx/36oSV4c+BMiOX+TD/RpKy3VHLktj4v
cJCUyTLwgIKfmLSa4YyRNfp5DlarLD0lejKJnVHGtQI9uFglxeYpaGxU34D+jwU/1KFnI3LfczMa
X2ThFx3Ho3Dp67PG30por5QVmcf3v4erUMwfn1PdbQ4Jjblo9FIR8XkTaGSCuoq/0sNKXd8KJtMC
Ttj6HuDhxUo54sXZKuPOmpE4gJSbXdddGn40rMSzpreMiKB9EDkWkOPl7YPAbfiQygizY3rsOQS6
5RGfEtIAME77fjdiPmowy5V6gEsonG1OEc6rT9oZdyj4ezDIazlJWexbDeipyrDi8k5jnutLGocm
5dTN1Vpmfu4HSWPOCK8rS0f2Nl4gqORfr4p5FTvzOCoTyPYyCjnIuOQqoGJeygdJUMVBb1wElyzB
MQzuuM0UQbT6x24OMzWUiSfW7w9UZnIwv/iHTzxzfgUh6nMmjohhu2HHaVg53666nVLG2HXcmfNe
5vBXtxmDEgEr2RB0QkIn/f3UrLOwhFsZ1CjYMgaxx8/OKAUHZcHDJFXHPzUu7p5HKQ+9ADvi4cLz
wgKgvK3n8ZVwUK1Nl5A0nUMCTomyZlyTIQP05A9zuf6ya3ED0wMJ8bmJEVxgoVXci6Q5Qy1Thjpf
lEsF79LOM0xJW+NuZ63YZGbdizb7oVPcznbYpVeroOZLOE/9FJmpzko+ajtvDBpC7QQDmXu4ZkZA
zUpllk55e/mxBEkBEQIP3lrUPcp5k5qae5L9y/cWJe4S2EMoPtvCAJKu7PLaDwSJGix9qNI00m/h
W/DLhzRBUQMxtxNEtJeuisCuC8lMDOGiXAg/XwPxgzD9De/p52PbjuQPXISZmXI+61YXF3SJ/eRs
5j+JLA7uiOtTkci0hpg3STRiQ0LF21GfXi/gbWNj9weFXmCX/MewbIdTHoEGqbG2RV+ZPQKYw5JM
FWhM9DOKD1w1WuF69RQT0FXTHmwAaD+ehJQo5toJr8bTTOWL6gcDv0aW6wdnDMEvC4us9tajuJs/
lGJMStHO7OKkjS1yyZrSJ6k/TaP96tdI7+zXz7gZBU4gAjJbZnu8lvgQRb+F0OdvN0906GmUdxi3
DQw1i7O0x8sAvKbOEtz4jKQSca+oIwhrZ4IPCQ+zScC7giYykBp5/3LBFf2Wm8fsjL8wa95BOBYw
QwRfYi0sJK3FnoLoDGSLemFB0JuL3yPFWTp8g+UZ7luFw32fIvO3G49WM9J9q5leUlnkZw6/TIZd
BMCy/b1oLDr/ugww7Ri2w9BA9ZrFpnBfR0ami2qBDjh0OHohvZCZ6fB+nAtM+I63Zpz/QVLP9l50
X2QinA2wQz+kWyzou0RT36BcdDWOs49BzAv9O2W2vYOiJE0Z13W2wv6raiYhV/YZFCH0VrE0p+t5
vou/RULI0P9lMGMgTy1DvERdIBJE/pyWr7mSQTHVUA5cNE2o8G1xv3G8A9YjUZRMeR1LstlPfkg1
tHUOc1l8L6GJfSgGNgR+oKRsEKVm62JN2KDsipacArJUntxOWK3+T+GV/uvM+3ph+EHznUEanqMO
d/rK6Es+v7+obPgr3JemnE+6fivdyZX1bYX7GnmaawA9qFfKFh7l0CuzmM/fk1mqPZth63knla0C
/mmnV7ICcJ/nxEm48p+PmzthcPjHCjI79sOiujpL9iaelssFZlz5ZHr2UyBT3kB7qd8o2cfUgBfP
jHfPDMvHXlxb9urNE6MPTevofXsdONU31vrB8emYrwtLcLL5G/gx8iBgFvai7DZHRFZkvJMwrRYL
FxDrXxAX7+vD8r+u7qLbz+YNAM1ceTVxYSm+wBPF2MmYa32QtcGrZ86+FZqdXxlY4CJW3EOQ6mmD
Wu0z4xFMI+MuHY6XcEtmeeAh2ckWRRI/lgCNsFLy4drc/eoOum8FnPV9vkP6yfRMvLabtewLsODw
Xmr0Zo3Q7H22dXNXJP31Am4Gq9nFsYTQpguUJlRwZBxwFIdrs1vKPugJGSt2Jrrdv6VP9uuKLGsj
ZPl2y9sEiMfZkTct7aRkI9QGnZ/N5q74ENgOzyIfSQz9DNFo6uhrDRSHbh2Ltggaaus7F1mKb3Ge
/XZa+WzV4SH8hE4X2PGt7hwEKDjx628+QHLx4P4HJ0ShMHt/cgIICDaqAX23LdrB+4WK5N62AH5f
gOzJoRten+bWWho8VxRPqRyrzqqv3LGYRlRti9NmmFXl9G59LyvYcy+f1NUigtEUZC/IlW9Siyd2
Vda8k+nb2t9Pl5VtQINkB4PYt1SoALXj3QJR4WDRQoIadsGRLKe7oqkuy/hXq4ShaexPGLydVDoK
dNRUldoJTzKHLAzPJpky7TyaKy99tAGhyxE50GPJoAHIfitqdJSQkt0E5zIPp/EkQ4btAz6Zaiaz
yPyrKO+LOzbcQJW7o+IYoLX6Q38GVI5snDlIKJO3vLZxKeXWOz0/CM+J7Iy5XIJByl0hEx+MG0+f
rnMv6rjqrOLNmR1T+1Zg3VxzSQ8DH9AmSEFx0HcTAApo5Z1S9DQSJR5bRAtBFd8H0+MYVfYXWysH
AFzHcQ3zdOBcRrsmtu2iSjBhQRJ5ZKjQQomlZCdD+FVd2C7KWYyniK9+xuKF7s6GSlSTtJyIza2U
kTTgvdJwokCOt05FSdB3d56yfpuFwXO2iUq+pKkrvvuShJy1A44UDdAM0TCTCfVPmePrDjX2YcTQ
cd2Nz/VoDDrxMTFUV+MI85OALyguKlGhIUclp06EIv8vW8sc9cnmPGMmcQm8Er8gzeeWcCScQHBu
qxJR2ilDbMPHdyrmfy10BZQDh+ZOmOEez7kZpRh1xWV0wyOgcPGcaVkq2e7QCNTv9CQywQ3864rf
3ekBCifH6aN9HACm/mkp9zUbBVPLCmGyf4blbwmPJP2StiLXRvXovAKRfrLVH85579rIEpDNvDpm
0At/RYArW8ruFFPt/JDIFzI/tMuktkdcfXzDdvqhsaHeLcT7EEeQIx4mcl7EGjz4jfOpcEy0Jy1O
e5NyhVeQ9WN5cUZOYhEToXvl3LvMmxFhMB8WmYBUqTtaISrmHeXVeO99qnVy0irhyPH1vyP2QV4T
bZZIrzobMGS4OgdN0Fby5Ysv8CTvk7xnlb1kUMYWtxwApQeKxpLmFTJNNP3MIF5WVTCYVD+/Hult
ydZT8duXDj3GaieO7+sZJYadMkt6TF3B/qngVQGotGFuJSX1nU3aKj2XiOBCAxVpj5PfbxnZ4w0b
su8LnXem2M0r+UouWP59ESQ7ngIUQLqoiP5aC8y2hxRQE3krWnoHRbcIPjWgZ6N7f8iOWaHpeFgx
Fb3N3A2BRRjU87bKgWiGfNeqNtbTRCZbg1XYnRSsMWi+nflUosnVMKYZHy8e53B3xlGs3IMc7Hce
+DU2PJikKyvIWLS/XYUFZu0EYsp0fmJurvh8NY9Hr8RzXfahQ4/+wnmrKy3MX125dr9ETW78+/SQ
iyAYTxMUXiQWErE57GQpR3ufWqDET7s/yf1yYU+0eiwIxRIdyVDoXizOdtP9LO/TQmWvyYf8dTl/
nfUZy14moQENJNG3/Lo7SH+dJEnuEIXD6VTtaITkuzpg4wIzuoPZTbOtfGC72fz9NQWNU/pQf/j6
EbbKDbGlSjj9wFRHTncX18szUjwaVhEfQfRMUTzwaDPW0mNMm4NX4dw6d6+bUt96n9aIvwqENL1Q
y9mBEmCrZjQQTO2kg64q6arw/zrjCbl8YKrZDc1NeulRe6rSLJA3RCOUL+Np8LDjVuxaxxBK5ycg
LojXnl+MLFxQzc8MgzwqwtuKEx5Ah2NaOa3Trf3D7N7+RSYOMQJIE0ArJwF2Pe2Ln5C5aqUVa/Ah
Btc4qjKiN1Szjih8xg+lXdhG13VaXkfLMZr6MlbJiTMKJuJN94G2KSQXNUAPHZKI8YYCAM2zbQwx
O0FfNO3wBV0T1hmAhPGWhXOz8fan/90z6nZbMHAuvHNKPrEbea2Dn6XqfEZ9NhlRWc3mbds6ccmB
GFpRyxFZpVAYw/tX1iYPDtf0KCQ0sImfJr+s9pMzj13xA1dKjozFCmlLjKm0CtToTMcRj4IB7OzP
YwL04z5F+RHgiyLymnwG9bRuvq+Z1VF5nmQVmHCvJmGQISYnVAljkjtTgQVcjpEz8TjT/eZXwkX8
fS3asIcyI403wxnP2fYNo0x923iKd/Nuipsie0XHbEPzD1s8Nz39hbbWr2ZIuHKUm7KUwi78UMrQ
jd3Y/+eOFqlDhKG6LomEPGofQBSPjRy60NLiLL+M8D6RukUAEVTxjBMCt+h3TPfrDJVatX2nSEpr
J3vibXoOTIYy2SgTDBSwVRQzA2vuyHUYK7QkaTgPn9S+SxAELkFuxzphDkBvS6V15XMrIbtWE1g9
V66zTG6Q8D8Bo7kbr1O6GZMO/D0tVmJ+WJTQ2iqDU0sVwlEyNUs7AuqVZotMLMPSv+L8iajC+UBX
W3gNaEP1NfGA7+rz/mInQF97w6twkjfScNp2yUUJhUTBC6dD4OaO8es0DmBhnC+eqfw6xX0panBZ
To2u0RdJ0Cjl3tIUraNCdFVVoRgsdrNr2sE/PjO9KtGr93RAyudHCYkAHacPp1znxSwvdMhV9ExV
tm4ONes4QTi7Ilb8Kyiq8e+FEt85gOSlDHNRhABILQ1Cm1bc2dtuh71dOKzho/dZtDCpd1r0BG6K
dtni7be901lP5vxli7gphdjngHDkWcKnbX7h71hobRSXh+NvasjZFcQlxBmOLw4sLKGXxc3pcLXq
QqD1vu6Br+AbqVlbW6fCd9b4TzbOm5QyopuGQi9SImrTZt9J58W7hppeNAy8O14W8HZB4PEeRCiT
TPIHmSHdF6DhArHA4qDjkNbRAVsa/eyXV+vsFVVCDzrkPpLyWrZtmVC7750tzkyYwYEYnd11ZpOj
9SAsT//VO5GRRTIp2HKo/43tVZr9Ob5SkfROKrE2gPCKf00mDoProkt5yomuDzlrt6EvSQik88Ar
Wt0VyjgfYmCx9cgr0qX5VwxLm6n9EPRH6OJnIvmEbtrZP+cDuQSORBFtI3KKBUFnkefwCu8C9D5d
8153ZH2v3dn+fWuW9xs1ViCDmR0fqdxTEnvNrlo7c9/4OkD57uphoKtfAJeaF0iJ7hT70kG93SoF
/7ENA1tD8K+vsoSaTTIMNtLVfTJbXY+7088oyAVdKT64lIgM991FwBJnvnatxGRg7DxTV35mfi5+
xdKWpv15sOzADmrylp0EUovXgbRfUyt5q3//OOSXn8zCZ8WudqdBXsvliX6iwY7XR/Ocx+TOOWP/
lBwlqmBpvUc7HPqdw9HJnGrYh//L9f+zAhIsu1/x6Xmb+qfmDaoR3Iv9b8PSewwQVUWt03qh6BjD
KrmzseFpyvW8PmME0MbeERbpMJEFp0Jep3sIprp3ot36dBNlbyv2THLNR/Zzc6JXXDQ6yAC0apOT
+xAKmvNwjNYgQMbJUqgPwhXOQ7CNHsAyw+n7OUSJXBXQ6Xg6AUXUK5OryNk7DRwE8eRxjqz2DX5i
SdqG1XBtqg8/6u1I+PSbNfwN5evmkgPWT9LSP2pGzO+RiNe2FOtBe9MFXqJKNk+zEZinUQs+7+Oq
DfnTjwlvoh/Md/78HC87VHhdntzXnEnFugKMJUWbNvaz4TnB8VbQJt1IPH6FzjLcb0dS8PzLvQhI
Dx9l6/V+wkhWQtqGYihg0std8ENRl9Xmf21pFyhgINY6mbohHd6UxtQF1FrBwFFxAKcLBXiq3iBT
C/qD8B/zKpj080Aw7X6RHl87AeO5xwo8tuP0xwHpuwFg8j0tDK5rVGRhciOOTHWvPgGDTh68/9j6
vJACPBnLSxb7mZCF8cVnmIecSjcnLheIWK8XBcV3bQKZGUMWvr2FzEtPb86GslQFP9js0HlcdSpH
wLi6qd5OgkvphLbK5JCwsm4l5l8ugR/D6ahy8l+aHVs9GfWP1ABAhcN8KGsymqVf9TMCwNMwOxag
Pw1moabte1+jWRDbEXZcoMtajg+feor9SvP6cpzFuTc8h//1927ex+TYNh66RxfD2L/kiRYkfZCz
O9BqnH0y+0pSa77petjm33RvWYrjx0fuTqvGEHed4ohrOC5CkBmMasxf6oMU/P3ehB2Y3HqL9MAL
qY42D2X/Ma6aKeNYfHjIkUENpw3OUwYsKcRC85KbxkFDsn2Zl8R4u5DvTQlDJ38TVI61y+R//SK+
0MVCI3/SgmKup9ApeT44mhDjE3BKOVyWHI12EgpYGajM2t15AMD9IkHasmpjMIweAORVmbeyfG5D
HeTKUfCbf8sOwHgyt7/t+F8FWhF/aRfAy3Qq9FTYjfF+89LY7xo6y59D4ImebLNKbJN8XqLRzwoP
dBiY8CgaRwLpgWwmV/WZr6WJ9JMp6YIZIS21NpG2gs9mcEMn6KBcpy/i2F4OovmfLntDy7oZ8hvk
0180YQo6sgky9R3b5d4JJf7FLFe3pp3bYprrN/a8TVdohjqM5v4Jz7a7sp6vmbf3ATByxzUmKKeB
szQlV+kHnHuz4hT2Zyee3KiUzoHcU82GnsQBzI3ShW+4KcdXyrw5XqM1Pmhr3NLsPAB9s9yUEPHr
82YKCETIZhmAlLvwny32hB8bNa91Y93xohFKYP6eqCSoiOOGRDUSLkNgTJ1HWWb43AuR4eQ52lOB
O9OMUpHGq+Y+3BbGCdVnP91irLao+veQW7bzFEFYPiOtX/QdRk4x0t8BwXwAdgiLyRLXC4w7Ym9b
Fm/Vtt2EuN9m9eA3Yp3l06oQv1jr4RXu8T/fHuX76oVhVC/1b000B/RUleLiMIWkR0T/2Ow0dlh4
UydY9rvEs/ef2aEOp7vn1ltNX6v9H1jrprUUhor1xDcjqNzkIG8Dkt6MToxKd36ZRXszQyHF8/ZL
TPYvJFADseIbOTrWG+60Z2B0egO1vvS36KsNTBfZ6J/n/qI9X+sXg4ZoITCIGgHg9HxBETgpox7+
zNno7AE2uJ1wVu0Di29zNN1yg8ueiVRZzKFFBUJvkrN5/Okia+OltT7gBrQBaTfIU7IXkMpe5r/c
Ib/SWI7e1MvM/8hAcR34eLeWop8mvxH9jFB4oukxm4AGqCRjA8Z9fao8OwcZzfa+whx18EKuHDeV
TTZvEKzjZRqnDhvr1mX9aYv0HtHcXxFSImkJQo8jXeJ6m4h7Cn0vYVMA8EgpK7u/++Y6SgCH1sE8
wLi/Xsbe/dXHaQe6J7mhaZshiO19xTUGp8LxfcXg1G3s8VWFpR+y3f1hSOWMSnVuVwGU3dC9V6+F
4OvIpi22+eNXD3rs+5rah5vokbtT11s4CbagJTkWIrP+QUSluL/pFix3SOUrl2Hm1xoLeJyHMOO0
IBU+mE1wC0/a+2swKDtGWQoIzeOmtLQFSC9RuNGzFXVfp5Uh7Ee4Oe/d9qHLpeS+WLbRwF5DXUqA
boweli45m8kKmhGtjzIFU5sLooPFPTJEuy+kEJtAayUT0e5a0plinaA7/hqqxpmJm7GkrNvwLrcg
mobeuoXknJbJ//5fq5M4ZbKJP8nZZOnGULyHygdqTm5Dy4nxwHLNGLtmvX9DaYjmjVWQfWc7+yE1
HWVgsxz4NBxryRoHTZx/ZcFqqwbPhl4TVSONAbPst+94OTODOhnys6GvYNNxKtckzD+RkxEjfVto
KpCHdL2+2H7r9L8ZXjn8Ev5NVjZ0/U11wrACO6qMzpUtCwgCVT543JTsvIxZOubG6TRD94nTf/S+
4cw97a+BY2agYw/v8AampDdT6E8bVczYPeZ8Bh5dJwWQdizfUMLDCemeLqm6YWpjigeXvUxOB6Wa
H2tLR7VFi5u1JyRsrsckbo/uiJ0yKn42Nt7z8OeJGu7jcCCZrAh7cUAILOR1/1HnnD2uihWvY8Zr
rCBN7VFxGO3/xRYMK5uhhFXv0aBHKTxLGx8j2cNtTI5SXgvGzsVA/po+bBcQXRit6eZG1/0mgizY
KHKY9XLdbOcWz1LE6GQtqXt82jnEk4fpjORZRzVjgHeXpAeHBgIExcUF34GzumXx3Y0o4SYhU6Jj
n5UZxs6R279+Eb/xQSCy6hQlOYWg7/t/Y98zd895XqjTqoqt4/yFT+zbQX4g/rLPnxOlUpXmEv5q
EDGeOBweir3a/8PsXMN9cD1VcBM5OqNU2pYBsfVRUTf/dO3Zkn6079jqi440CfEG9TYg+qdy6qds
4xZdTOPyBa6SQPRWzqvV0ljXXj06L96yFkmicvzyobPGeR8NSBYW+jeQfvaU8ccpT2+n6VIrguWR
sedDKQ8YqfnIqYOI61oselziwQVhmJPAZu5NCdnS7BM2/dfIe6Wgn69MybYVZZO5Ior4VfzI1kEI
+igbGBSFdvaZ3UOqPXVX87bDKwAbQVt7uS7EyWkiAq6+kjV4xhIUu7tRkFQxW2GWEwXd4nmsRZWN
fDJ6Bu3epJL7aP5s+m4YA7klK0TPelghRjyK0KDpqoU+pZxvWWW49MqNOlsxwdBokcV7XXzkJZcI
kJ4uHUcegRiQZvkG4jvDjQ+Q8M5YbQ6KsWZiEp53T9wS3eDQa09vsPIV724DioxdCsut3zbR/ld5
iNWid2u0rxo8E/E7O5B3uRu7M8+ihIFXdMOIzUU2o3SyoP1pd4pOlOpJRuxjTzizKum7DL43VjEB
QEuVzOOvKGRWwSXkW84GwQE5nJvYxIIbKonO2qRscw7JX9UyhDLocrqupsAUNVp7jYSissrLuO3f
PqpZtzBhDus2lfh0e0SD7BihWpKECa7XXWFaZEtALHRLY2L3FUZhkw5IWlR1GCt64b9XQokkX1q8
RHSUhfHxxkeQogV6gQBd79TgGSSBRvgXSirmn8AyivBHNNLMk6/MngBP5D9X4Ktcug2iF3Ffbg9b
DxAX9169I8HQERjEXSpK574cTbSQ+NP+9azpe+HxqXTiS+o8vTj8hYNG/Bfc4wV0jI2uH0wBh3Hm
/OHyYG9AFVUbThlhEs0l4gaDw7Bx40X1z+/caIf5E0pWskD0DtH2d82UxPooT9wc7U3bicGgmVAn
sOEHER4XfvcnOMskYPVGWJiX3zAw3h21dFDO9z2/g9cU+Z+z/0I0R17R5xDJyeFffBjeT34AdVkO
YYDQUTVF1jO2MM8H7FIeg/5qbSMGiY4+sDVzwhZQ/aswTQjaLpFONYR/E6K0uUNhV476kykYWrR9
RhQ9NRNHkzcCj/ZTZE87MLACti2EsvGJnxo4dupxg17Arp4CzHMnYFJlgD6v+tjxp6C+VXUvWPUe
o1p03hw5NHfH2L52kz1KrfiREbSbiTjbpilYGnkC7JX50aSj7PlfGRZ+RCEHqgeWfD3QDf7pbGA7
tg7IBblSo/goFdsHFteY8jB5bfMebf0WP6crsnCFUTG+YnloALQRlBwGnFDFf+WY1ivvjytkhjsg
KmraqfZ9yWAM0lG9ykTiARatpEaAWdsELQCmJ0WksgMz8CHn2iZPBaVRDDnfQ6RSHz4xgsrmMz1s
KEyPGFj3bpE/BSbpAdAv8bdTelLwv5WhVquVeOkM/wUrtk+f2IOOW8Fi4Esn1IEGeHh2toKMv7s8
CbVwb64hNGoJHA5qrr9xwgInyIktNT9BU+u4aRs/ApEuMop0aOXZDsaKvCEKzJL5nVO7a8eM3AKW
SP2wyvlET0LmPViWi4hxRLPtfBfxggMRyfUMhGeVu5Gp6qBkt8f2TB3RHC3TZnplGp4jvvjdIC+s
8LSNMnlUbbafOmb2mN9620UQFIV7HtQlNoerc645RF4GabrDcE25RG3udZFN8PHMdm8H83y7oWh3
UFUihgSy7BdvStrfDJJY9pd13mLobppWWf/1EfjTZ7IgHR0BuB3fJJEIk/8KWlEVdI1XLT7Wl2k+
selOLvp2xd2XvZYRsbxPfRhaVK+3VR9FaIwG2gC0oJgD7VBGwPXJh+7BAYFuV2ProhroBGkKRP/y
DOeOa0PR/VK/de9U913DiO+3utDCtVxZ3Ab4NT8MqnUosv3PGh5P6wZNaIo5oCqtRIUMppS0B5sG
1gU1V/lWZYCboVLkm3LjlqqFO2Mf6H/JN531fPzOrte9LgsPKSMwE2nXpxNpyt1+4NqJb1vZyobQ
YrxJMoN6WcW1xpkRTYYgQSXZMveINhrLgkDV1l3FJ/6+aP6JT7axeAXSJfgsZbKmk8nboJM+thFb
xJpl5d80dHcH7RQL22/q4cOkERuaH6IamovpUifbY4c1VKEIdHEmTU2NXbachAlRTZoBx0cMoKN1
PCOdh2xl4wqJixiJyuynz5IF79XI0err9obHXFxpEPQclx6dum7fdbQ9ri/uOxPlvWfdKOzTzDOl
DftpATqvOknVP61sYS8AX4uIFS4zvQ9MeXqkl1MVqMNjxg6UYh1WBOqC16IWtUpsNQK3DIVfLu/S
nQIlw330cxwYv9oHP+uGaHG+7caeSqZhpnE5919/EV2REpX1Wlqyf7LOb2YmsEQWozNqCwdc//Kj
lr9sI8N4+whCHNz2r/PaaxtJjYrw+dUx3The8WYWqlVMXNQ5CufHaZjbKlL2L+7CJ+IlDLKOWjvz
pZ/JHvLDtI9MQ7CRoDZxoARR0cwsjggPD7+9ZBr9LmW3Sb/K56Bw3FvuwX0WIAlL6Ea6CUh4Sne9
wx7E7S5I2cPQGtbz5BU29Y1yjij8F3XikjhUBRjCcBeb8KVPnNgywHSIsk6hOO75NC86cqor9PTK
6XVurCgDL3yftz5xMyfWQpyZY+SqjqsAl434V/0hrvOhx5HF+y8jFMU53dkI32Z2EE3cUGs7EDLR
3tV2kvnyYKjww/tje5bzWYxz2cIjnIq1syGi3Oj89RdSkVxyVwUQWr04KnhISCnKjvmDtrD6i9Kk
TvaAkbYqLILFPsicc1kSqk3lNVnuW0xeYsBTBTQTdXvki9uCquS+ds1xdIwW9nw/lBS7QX6eoiAj
8mX09biLShi2zBGqgg6+3BQnC3Utw2P2IlGctsbiQRcPcRz3yhRjezrVRHz2Fal7mX6oZGPB7tfA
DuNQH4BT+BKg8x2wsUMw4EyQVSRFgq8dWsPnqrfgUi14TDdyiPkQeYvBeUslVVbN5T6N0jpsIKpN
ZYfLLVTlpZnqKcy6kwa7mjKW2DW1d8Rf6V5vSoWaVgRV9uUbd/n8p1rGZ0DguC2XLHfJt0E3ErxW
KyRtC2iK2Lx5p95j6c0ABCu7Ob5uQZLo8j4VKImjlbG30OTC0uI1Sri4ftoYG6TTIkM72nHmZ6as
5P4PwGztRyuCSHIjYF8J/ArW7j+fZOxeZLcxPr2NGfAFwYbnyXZ5gDgGwG8Vgf6Y5cA2E2bosugn
WAqtRA/VMSjPw3PCfntxDPgD3r1495A8GL0sSYK3hGBeXPEIF8fa5Mj8JTl26W6ESti4RQ4VnfMR
hH6zU6Jo/uXw/ZKJ3ps5o2rfgZy/gPWLtUV6T7idftLJQkVZa/anwN1LXU1MKp2C+G3u+cRR7Y6Z
+2pyssC2+Y/y7fZBNTUNM0knVYX0/lTn4+QZuGWlXFtuAB9KHsTOrCz1tCINbe4PPHC6Oy0urWle
WnVDF7sxX3sRN6r0WZCa3qoCJrOKHNXFYWrV3E46MwwAIZVQ77yp+vIdapG/lLUfgv6Fb+SYQke3
gnMhp9FlTFeDDii8AoF5a5bGDQb1NTEYAIQpploxbod/NPze3sHUJeC2XIgRXv00yBi3nrIxMrOQ
mUFOObqgZxsVWD+1BFD8VZ79WEczAaYcOLs3OIO6iwMpaaujeBU5f5eF/UmYo7Zx/SsDHZmChi8k
JVuXIJjlG5CDhbcLozSUmbq3e+vCuu4qg1OKJpz4Ie4gukDUy0Yq3rIB6Fx1v/YyvJse1u1lmqhw
IZgiQXMWBHreEGC1Xj3p+0SMRTrvVjh8Buyk1gAj06DG5lDbYceCkiiwdtd8RMxZPioXz5RUpsWL
o4Rno9UumVr7+Z5ijl3WsopiBevWtXbNdfl7y6Xaju7XxuFY9mxP90cVNr1sCWZvCYxgRI+a30z6
5nc6Vh4CsMsrkwMieC5lddY5tXAiU2q+QT8oymiOdRp/EDoIilxZufzaQNxLkSq8PFRphyq0Lkc4
WVwbvSnuNpi8FzUF0dawnYkfmTsikjja9Hbrpk6gHSc5XZqE/qcthT7hS+0b3lZYsamnKER91aR0
MnCkr9g7E4ECg5/HTPTpOkSRxe92vryAe/2W2NzVi0n8pMMg9tmEQJt37jgn2j95aq740DNb7VzS
eTcQQVj6jAxueOFb5gc9XDOydzcwtiMPI7aOPx4s99Qk6Z6/GdH1qeVZbXIeafmCcE1HTHkTXTvF
7jUwpN3vXhIcuEz4I3Y+XqGIRndfuA4xPZoH3ByxIQBYTR/IB5kSm3uposD9ShRcni70dBlXZYBK
ZsMCOgykVeJS9qNb3ahyEwBxt7hSmBDkDxAEuzodq3duLhIr2fwYYibjKsgpDKGJ+QEiG+eKxJ3F
/D9z0hAA+l4Ch6txWDtZwu2HRJzgsiTizTsomEwhhJ50c8UGIDK0hbpE6tBL7gLulAK9HwyrPS0m
k8tJd9gaoRBHQrrVEdle8wpye2HwGfXM2sRyE1ge2FaMhUra5w9ioYchtLfqTgqqRq6p8ldjRKOA
UT+n5+xdWpRNKjkN/Vnpevbpl2NmFyYx6pMiU7icEtkbA6OjitHE7EyAkoQeAablQ2beJIZ5NEZ7
CST2UN1I6oEMMmgpBa35qiY4lLs/6QwBcsB7M2VyDsRFsqYRmFas4CKyezwO1As1ehpcQFyaZS/y
iB2GXHxSx8hZLkq18kMuc4Ugyw+rwYqnGl7uwKs3lBuTi21SiLxbaVYgluPAJ/K3FsTgke6evdoz
SSpMWPDGk3rjpdkGBoPiftrVVySIlyP2Ypdy/vgzwzJa76ebgwby43Z3RBNNeI+vVFlHEhG8g4ET
C3/qcdITF7bwxdhhLsPdFvBYyt+IQMoOJ/LgUFqoDb04zRcF/zT+0NVyYY6mgLMU3BetVM5rCBWV
VefdMtfabW2ckreGsVcW21vWO4FV41U+LXH5EeeUHZrsEfNFpSamMwOGBWdnWYa06bkn7KPozSrj
SywUwc9KzMhEFk2wBa6vS5VHvTMhf6Jvsp5103jQHmX6DM2ELlxAsh0YLUMW96sby1wD0JjZaEpi
PGVYTri642ACqA9NW0ZM1IrgrkbKtOzKwi3CYLsqYTCoTi4lfueDCNSmFk1WYBbp9mjUnye/vrt5
FhwVRnqm8qhzEkyv7ikf0P2B2bPO9G10FqiqXT83MqzajdemXfqY8yLSFKIh356YvIaHvP7Cso1Z
OovwCRBafskCkCVcVYf2Jf4UexrR44uWe0cALSGZTKv0lY7xaq/lOUQ6Ynm62kqoz8xdJR2r7lXi
CkNjqRSpiGmHeDLoIjRUJ00JYTvt3/A4G+jlqeCgILF14/Zo0ljaZ97ZKn/jhKFLydN2hQd480Ur
D1AbsoKl6yW3iFuyzIaIduNN1lzfdeB3hXa+Ai5JJmUq7vDK5zlStTLtDsF97Xf0kMrne61cc/4q
Ll5SSqo4G/OeyrgJ7KV4/0bsjj2JMGzY6Pk0f90g4RElmeJAShV0lpqGYXtpuycPOH/8SSeGVqSz
WGaJexlqfTH/V/lgnHyLp73Yyc/x20RnCxLNiMoDC8kfZb16IDKdPPN+6sG4hw41nwLZZPFIX32b
TuZTxq4rqdp5LRAvWAfqsMHiebcrRAJuXoDmclGPCBb+wkAeRY+PfCMpf04GzerGi3pLN9lAuV3D
c8wRzcVPV7GkcPNUyQ2VkDu6rtPaBOjGZAYUhbNENScGOAqo6pxtHCU8HJQ+fESjuVY7bcTEXkq6
o5fHVld9iotYzRo7DpZAB2GTkOpunE/7rRLnkm2K2w+rEuUBv9UczWBOELCgqaJCt1Jy80J+Fpr8
bmuwSXvOjeUg4QpCb5Dv8qfHoXdeHUN44vwp5t0Ik024naxceRQ1KCmpTyOmQUgRM2vZW82CgUjp
Zo9Wh63F9rvXjIuKI8zjktYNi5O4/4EC/LNCRikZr3uu2xNGJSru2FyGHOiQxrWGXoTaU1y6fk+7
0CxWTmB6QTSCLMwdt8Q/x9DYnxFbhA6kfx9AimT4F9Rgp4ukO5vZq+PQvy1we8McVxywwfz9ozQs
hKPaA14yWLYhpyO5WSiFjzD75DikSSbwSqRsL5yk/+gk/LR07DMOgT6dvwyVdfRS1uon/eKj/yPF
wl2sCAkm6hNJ5z2mNblbFzULrTXuNDIUPvQWpHDRrTPgxysfZQ7PA/50ini0AdrmPeTFJak7kDlM
o5FQ9SqNTV/7iP/Uogg5zkr1tCWN4fBIrEDlI/GR7S7hUiH5CMGPU3rfNaFRy9Vw06JYYIxnVbSq
ajxB1f9wPWTlDushDSrFpeuBt3MLgzVvzgDXM9VELrgY2t4a+0rrvv/i7dzc8fr4+MMErgDBrTid
N2Pbz05QxQ7HRIawJb0qUuqF+A/CKhD8HoOU02ABVgp/DAApxzhhUWvjAaIsl0yyK9pnLdsnChMK
VtAjntdi4Oq25b4pfwBK/FEZsRA97teM6dk0bc88kJUPlq9S+h9emFS1BoclRsSix1Rh6vuM27IY
Zw424HVe6NXixZrX7qoLBEAXC2dKg4/oFCAuwd3/LXTlmM0WKT3zV7JRx+D1/lPXp/O76IMb2yld
CCJQtSMkG7Mcu8WQNXiIIV+Fut6wuu/9oROXsRHk0xZFeIfuFIgKjYS9+qRfryVMZ+EUL0KgXzDV
Tjg7tH7AKwkOTXkxCLAsXK74cMjlsq55Wywxq9+/aToTM4DsLVZgr8WrlpOQTlLezXaJYRXWXwd+
/ErNSbCQVcC9IeyoHwsOqRkfCRirwYqY0J+77NClG3AAal/iDEoO7Dqtctiwvhq47yHSEA3sgSuH
KQ228IUdd/Jvi5IpPPH3CoUwuOVohW105t6wEI3FXSgfvwN1gyBgqiuJ4jSaut8nMwD0UVvOhWl+
XnXMZaJRUz/IpEKkTEAc44/xOpY7oUFfCJhwTBk9OW1Wzjmj+dWLVhERqS3xT0um9H4sg6q/d2+R
reE1dlcZF170LB11CR4imNlYt6Ml128HN1AQCuX2WCXO4Tw4rSaHMT0DUvkZXoaE+3pYm/fyW77r
L6Vfl7BsZb7A8kAaEqBX6Phl9bjCIf+vRl4EaaS3MytXrAUtpDuwXjNhfjnqUu5SE44+Js/KNYZ8
ZSnOG74vTntz1v6PYMi0jFqncdRzMn4u5VPU7gGQzNGA/q5lUPuFs8BKgDWGjyztikaU2mNCSv6B
7Utmgl7O6hSvVbjuRErfW+lXmUfPJJZplubiE4DdU067PCRFOt/44I1xaK0jmNGQGvWhuN0TKbyW
hVIlTh3IrMj76+icfN7vlgN/N2MYUfTTPLvdhlpiWu00tjn4R/JBBGSnIi9TNBCGEAPrZPpUD4WO
2+qNJshwyUKFwz+LWP7geTprgEyC9vwfcFBK3joeQZleTm9gO8PrAhbyXn/Pgfxfq5yKcVTEutuj
Z2xS65CoyNHKfdcfuWoKI168TY6fM0XbB6RuY2JwsFUz7jRC4TMswM26NYLHU/9tbBVOee5d1tM/
95J3K+Eq2UojLj9qaPm2NQsY/2e9pL1Hzlyl0RrqU3NFBgFW9aFpanMLpxnnR9oYmQX0ZFzakJHj
rfmCO9Pb5lQBSrpJfu9QRC8VrO+iBg3vD4X3SY2HXPaxqgAlKeyoFw3ZA0WCF4ddp13S8N8WQGNF
FIs3rcVc/HWXyGQFyZfzETe1v28wRuSrawsM5wrs8UhkARbvacDph2okI5Tklam7/zOrgIktKHrd
hLEEEWX3a0lwfoItUFHCDxp7E0mlh9NxCEEI6bMrQX/luueDjNI5PpTOH3lZncQuDrKKoYOH8GKC
vEJ5s2tQ7Inna7ZOLps76mujbRB/Vreu91Tbl+msbmsDv51AV9H6I43dE3+m0iG9o8OlyEWh64g+
w+GS6cKWZuxcyBaGwMEHXn3yGQmfZW3GDw5wGTztjnOZGL18qeVt/OJXSfSGl+L90OJ68pKw8brj
VtHohLx+2SRmzuSwll8XM0D5tggZfx1Luvor2yu+QXY4yQBoMzd0qx2NAUh7Tx5uiPV3lcHwFZ3Y
UanAxlDhe2+fr9p8e9/MU1z6bIxyIOAs50UkE3Xy4zBXMAT2EaWHs6yTBbuA0i/rUTDkaqFBBkH1
X8rxyatUaahbvikvsJlApXS3iPQjhxxbmAO2kFpGhmLThlXerd4dBAbEEuTKNAr5ksQjfG0lGolZ
bDDzgWlLGqCtHT1izd+n8YHiZuOLGRRooRM7fef/Y1qlNbc87Ol7ZV//c02uvU33Xm9+oJ0wBiiN
UcWvAHjxsBo0RZ/J9E5D3gAeHYyfVu0yZpjhlmdIvSPk2jBHTbHHcXFD7rkC/wSAIy0dq/2JJSCd
/Acq6NgmOlubzOlVc5ErzbY7VBzakrxx+6riGAzqUEFsgOyMSaXkiMxA/Is/vJFlIJp1Ql6INhZ3
cJd85gbbvURM6cYLNaIanRwwwLOPvkbx2gv+P/ghiCt+vaeIndK23WlASmNBkr/L1e2d/uDHt0fZ
BPR22oJ2Xdot5+xPBGetwVAXmKSyuVKJLdilDhQyQWjmr3xxpQohCivs6YK2X4kkZL6UoDZ2sb7A
eVr/kGrmW3Ci7jfzyxEeTfR+YLmYMsGCRcv4x4eY7GlSn9RA6F7eJItnA7SjqeYUf6gdyKQDIcuk
yr67UAsqfKMx6G8sMM8ZUNrSmRzkBqPuacb/4lc2+CrwxfOaDwN4sFKOjcyJakFFHmeiXc3V9zoM
4i2shVVbwVaFwhxhrT2ld4HpUXTJS1PUSbiBbH13HdIdavpQTfOR31Hjqnn42t/cM5LnLUtDR/fR
BxpA8EpOfxYAwuScE9HJP7WVXcGGcM+znAThL+w7MNAXDlpdMqnqJY6MrMv6H04EcvbMRR8rXqD6
jpy7Yo4ttmVFGv4K29rAw9j/IhZ6HHRQ0duF0Y3SI7XF8Nppc164qTB7+DYOJRwd9Q1dDoeFjOTx
1H63tyfrT4kzcyzAXyPApcQYkwnrhFPSzIiqoOqaw6HZ84tIlcFsES/R8gTK/cs9ZcPGjUHp30bg
vuVpakcHJ2tJ3E2HVQkw8xUwJmfSCymaJ0NaDXt/SXnyjdtFeO82oC0JGFwOFete4GErRm9+w0NS
vP18RxeXJQ4UrDNRs72OBrIDod13PL0iJb7WCvg5pAZb+pMSnMKWhyfs4g8/8V2pgAIa0NQy4U9b
2Vqn5BFRZLQ8Xg9xwGJgZKi4r+aMVsYWOThKmTzBpRSj77FXxeOPCmRJtM4VEI5PWgL85rBL7ETO
sG9UowrwFSBNLIsSKMNQclaDb8+6j0ly6a6dM6/ctbrkX6AfDHBpwaxkcE5qDVEwqAYXhpR4oc1m
uTlpYYzgHPcw6GFjma4lFuU6KJbQ/mv2xGdpNM9+aMNQOAVpGMH5/dSFJiQgf9vbvbJKYhMtS6Y4
uZlTrI51jdx3KoK3gnrkEokwmeZJRM5kaf2a0og1jkdCQrg38MMfanY6eNnO9gg6N0h5WfMDsQxV
LyqDZ2MH5opFvEmk+2uaA0MEycNcM20CxHKFBg7C9LLdyUe1yg1H7cS3hxyFVUqBAJWs3CWUKIdn
pcToh49pigEIQwIK+kuzvGIjRwFjBTGXUmZnbbtwegT5GE5zsSPNrWU+tbNvrRA4iFai3+B1UKt4
ql0A6RZMuHHig6/bl7UjcqKqE7lXgxx0GULWftxeQ1IdczzJ5CChLW3tV47rcvGNCIDWc1P8vpBH
TQepsi9IqG4XTXZpPAMyaZPXLqGrTCDbfppjvmsppBLlaswEovRfGmM6cyv0ktsZM6s6boy6wZqY
UdIMTAvTq+bPhxcsH1NQ12gtj1Ky64RQqc1rTTnuVFela6RZufcZUrKFCxVHI6TqYA/GY2vAfWFc
CNp7aGQNBNmyIi5WkAjzZ238SisDtJ5Zi0jJTwqGhaHq2ztBciKRwlv3aVLHvPsQeg7rqRNHpFrQ
1dH62u1tHqsvrq9+yZ4pUQlJ/HVjemuTkSzp6mkxjYkngMioJCsndR6iElmzYbF3nqveU4qCrXys
39HlV1W6NdeE1EgbiGYNyC29ibCNKhkcaOlbwAQY1HdAH22W+o2/0kjyf63/gWeZXzOqWbnLOr5i
gdTkO8rqgOOVD5VtMaMT1+QMraq5drOP/U6B6NvPa3QfBISjSbMRI+LBHDLGl1aF/C4tTCMolgck
3uansYDZxzbdndQw8aoZixDjGZE+iVUtBiYZ34g4nIFf8nlO3XaEvBknof2THKOadMlKSOFNUwVs
X2rrJBz/MK/kUffxWdib51A7r+CMlGbieZWJw11g7FOZU3EztI6x5YZXmjHqvVADiNa2bW8GVIzM
4e/s37tGnadaJ2n3KIc7C1NoXo/jFDDmlww91U2AMDvcu2eSL5SZJBrjGN5YSpRbrLPwAVX95gug
W5ajoWgR6lhTfgl7Vo+hpAG5Zao/nxvmgDsr6lDWHa1vPw5MPkA7HpiGNa6ZP/+uDLyFUGOas2Ts
ekoxxbnDapRY8f/gquYhLvtZ4TNEH0wsNx6Nxi4ovcmtWgQ30fP8WPHYBUTYlRvyIXmigjDI0O3/
vRW5RGroZsiD8KtykruN4suuWueFarMibNRYrYQ1qx3wrRS5yk7YEgVmS5XR9sDTZiV3sd3rAA/N
0kQCThiulYaBo4OVBWx1EIgHHN64Ch+HDVM/cI39mHXy88BBm9uzFud9mUXuunIa9Ejfufx4986E
YzdeiJN62hRmnBiGaGoNSvSlLO4mhFH0FEXzziXdONc0DzAYv0gz+9oTGnJvPYzvSBoq9MsxPwd2
WyRcpst/YGtNfWxHKYzSICTKfdHVu/lBGdJFixBNYTFZhWFBWRPQiEigUtiM6MMw2IniGVQ6nkfj
cVxB0JmuHULAJRQmFPSi+xY6RsWj/nKSV1MxLtHNCZuUbg1iRZwWp42ue01ncl18K99lbjkswW0t
41iYQfvTqxD/7iO12Jy7N7drYCSLB83MUqbIxZge2dd1rwbPBmz1T6EHDDr15Z12T3PC34DB+mmz
+f/EQu4aQhrHwm7kMsu+mNTQJ00Z6+2Dba/lMUe+U5TX6DYsme74FQ6xdRDgmSWyI3ADoDiV6HEN
R2ALTwuQgeyxFf46MhYhrrlpWQsCHLLCjuRVHF+OK/tVnUQAeEtW4UGRZDtq9ZAy7SHCew798QEn
QRaO0Aqaqy1WJmNlWldXUKvNaNrWf4ey2yXe3obqKcFQO/GfMWLZ+VhdL6r1jGm/4MjV4UvreEPc
Advgfy7T36a/jXW6jl4bKxSnu1OkObohG2LtdlCPGQI/3AS3VkcGfgj8qk03PF/4oU6Ro7z1dvX7
YJwuWU4Rm/RctdlcMwaoTdyH8z2BMyrvvHOsQ15VqHrnvVtD0GWRvg6/Qu/hzx74iIhkMuMst6jk
THAGbo36Wy6gE3ay2INVAqSW/PzlDoESKL3KXwiJmB4LfaSg5xASGPeHFODSOSNnXywBOkX2MHkx
WskHn0qim/JTRBLhL+/BOXZ8n9JeQPD2D6Mzz2IUz2+SmSTpRCXIjN2FA49PjRhF0S+8+XSU3+fg
9N+/lFn1hwFkoFcyTDSgnC4YBhbrCESIUcjkAz3jheRytY+cTCB5bAmhRAKE+0ZTFbkQggQK4Yxk
NtPlnyUw3+BoxMxkAyBtHDZJsL7Axm1dGgR2UR8S4Lyttwfn6OUrMkRSMFTv9F95DSX1wzuklYRO
aoGEojWB9R/bVXgFHe7rYDIf5+cNO5IND0QrbzJOpSVY/ZS8Jr2+JH6tqLEHeHKzcS8/yUIRGqzA
e50uVT6KODPj5KfgzJv3dBUm+ExoZTmfNBYrFx7fxYRDi26hUKhD94JmZElGypmcFNMZ9e5rp8oy
ICo47xiQethdxz06v3mEfpG8AVabIodPJOAFS1nmAD/bai/DGZhzz/8+tA04sKq3UEDvOVWYxFi5
lm3PquGzbo4/CFoV/tYjJoA+7RryLsQLzlygBZ3dPTdJ4kF+3tw72vZSaTUhPa/E9Ia3lT5G+zF1
/fZ2po66YzF/7z/NKI8AD7QKmPcRGAAoTJ2NJ6NzIh/MrkJJrPrpMoZ1hCzhHza/09j+T5HByEX9
wPz85W/T3xNBjaFvQ9DMdYbIeMhQBwI7/Ahkv/YuW+B3ntMAE45fgWx5wYdv2VsJXlcHtYk5ypG5
OAK0v5QgFdSXVuWaWCliao4GEptL5ULby1hZCt4BIMiMpjuddsenNj3tJLmNReRe+qU1R86WAM+7
bnuNSM2lYvLDuB5mP3ZGbNdakA7m+bZZWC27d9HRFkd79x1AuQjv7HMAmp1gBvVyi5VEm/iGmt1K
gSFElNm0atNkj3hOXmwuyIyP9AgFrwzLvYbG2F1z0kIBc6WOeLEhGU5EYlqclINyVtsSr0RDqS6P
mmLahpsm1tS+7zI39KRledVxnTyo2beHiLi6xpIDY5au8oauaFL0Zdl017sYIX6b+p3i4J8R0tkK
tSMlWY6gGVhPCnR0lkZ7bBSFV0+7NvVIR8Z/SGCLtXg0QSsHEo5PvRjG6tOaFuVAw5pYvF+vGSCN
EDLiM3uuebOuy/MIK8RGV71CDuXn0ESsZTjZntsYX5CFbARhz+durqgAiBkIL6+YgUkb8J4DsWC/
2AlVMj7MMJamC4ukDbplSbFsiEWRtAOLIimGxIB3w3sG8Rz5YaTiKMTo7dWTtxM7pa5zsuZ3aRfJ
5PAJw8ENTo/gz8kQnZKjWbyv1bHhYaGKl+da7KXH9Ns0XewPAZMLS+z/vw8ZSUk6BEQB3wpX49U0
Q0GxwkVeKmG8RT17+MciHx0eIWpIcpJbZ8kd4vYDLy3Jws9U3Ctboc1bmwZp0CAA35JVwzjQ9Lnt
XoTTxqkBACsFhDEWjVBTZTxeDe09w6Nkdmgd8ZbfrKec5PuWAELRJn5b6GLPzYq+4VrVXmz/I6CB
XrwCb7GdWD2fW1r/sm72fXAyirEbKzxROEcJf6tdWnVS78Bp1K8nKv1iZAb081EXgWcJrIhGyap9
qtBckuC8/Ax0JG4yj5cGyTKRx6X0rbRUhBHvsvhHziLZdsD/dpT+sQ5FLpQoEwSKAquhXZZeItTd
i0b40qwzDc5TbwaCZ0Z52O6Hn0wpUcNupHkjfNEokC1xFRB9LVcOxbyYL7eN8Ay5YtFBRfJAAKYN
68lhLAkLQaHHsDG4OF40I5e1laEZhmJSCUbzOuaDse5PYf9WIbIlp/DHIWF7MM0TZ2B5G+UHTFGB
E5c+2BALsQlBmIZUOavlHOn/HpA9qcVnnY6CJCMRtIWSQNlzaGV8Bku9kmgvHpk2oBLl6GRIqPD7
tWWQ3wEY1Xcdx1jTfqe9K+thaKTzwZ3/ZlM3rrr/kE7vUWGYJr86uHpqh5ZeKZ+nQpdci0lmmiFl
qIgk8iVHPR0shtcg/eb58GhJoNheQI/1jRYt+LM87urnAJnHESwCmpZKQs0VE5ZpCdWFc+myIqmX
fawCfdZERJi0uoC4YUvfd9tmyw8/UM1fwOjzKYOUUzspx9XMi2uoyI3pp9GvmSiLPo/GapwsuMUz
dX+L0xJzhz61NcLF3/sMrcLFEbuIcELiJ7+dmRllT9rSQZagztyPi4F3bY14o3D/tfgMBP2JxSP4
dTB+iU/3Zn+mpmzaGunp4NwjYdLonSLsTLqexUlbgvltk/8eONsPwLKV6mG1l7Sp2pPvTWy25Q1A
AzxytDS/3AZqMQmzbmzoFiPpprClvaP7XLJ9Y9kpvwTiaBU0JoBajprMGWbcesvp2AjOi1e+pLLa
ZJQO1SlzRFc1N8KZEky5FOUt5pv7BWqtNI2yOtEBCMcEFJF+LUqvrHJ2tI/IU6DpQgT5Q1Xo/RXS
M3CWacCVee7KNHVa+j0ptc0eRawGDgFZjSv63UqF34WeQHElSJPWr5gw/xr8/y4mQl523umdTsKy
mS1QHEYXCcvHWjFSI4ycENFKsf1XTcGrUKIOyHQDlnSiL72I+pMtm02hK5OgZrbVNHkd40VeDdxY
bACPb0f5Dena94zB2YkBWxVojJdJERGyclJLG+upApg6hRc4A5d92ZSHSuOW02WpNq1fgHz1A/yY
cxkD4CKiJ2ZNw9LnaSnBPRGNuhglx3hAXz6Lh5NO925bDv/MogdXplmk1YtYWBkzKZcByOJmds3K
sq140zx65TEzR4iZQb1BPwcWChitFH6NcXQrdqD5vwlYnPGw1/Feu0Zd4jbsIuDMJIt8GJnb2bxI
EuxoNuwLiBJGdz5GY3wDRDP+pFassFTn6s5RONGApPt7TcPqu1eWPevKtfXCLKILCTJg0P7OGmlS
xYEKbKpYGfNBXw2s27wJfseCiOkmXewxLA3dgNbN+U5kMUVJXQrlelhvVEGSRePplwzEKj42wABv
7L4M9Me2Vhuo9kam0CRzhLG/iLHRRsQ3fgqwMygf461e7+I8PmT+OqE5zIakacduwFka3kIxpXG4
udJ1O3nebVfbPcPR7yg6BItDIo9azuhGx63boOs1EGkBxZq8acOe6MkpdqK4W5hAkuUWXDJ/x5Mk
Z9qEEEoxf+YzId2iWy2SbrIBKBm05BBTTJ9EEm87qVBs1lHz2lP7QzhgGauuEJASN07kO3ZIWkLY
vc8+huTER1FIST0308BMYFQ4mRpTA8PULwpnDQmm+U9Fj8MB8oFxXzM6WiI1F80MGXtex1EbLO1l
ku78U3AbA/oVVDIKoFey/1J3qp80lHMgw5KklDIABsZV82SnkLDrODxgH72MxZzjSW9BEtnA9LY1
ppUV8m0VVkbMtdV2XcPDxtvbbgXQ/Sr1cfmuJcPo8HEB/Oc7SeU491yBMWQBnLeF+ands2SPBhMZ
ImxQDnXed6UglqiTYYUafqQGaezTVIoqsGYgYuwVvkkBjTYAKHgAYkq9bMHN6httChP8xUFnww4b
HcdrYdOHEx66rjxfrUQbj+M1Wgi8UhTuRkiBEqFy/vltArMn/JaFJyYs2TYCsaXIsxk8oHCp10vZ
8LhV1bFKfvVL3wahzmxBwX+wpcWh/qaCikk/dHBcAKO6K+boD0qK6/aqBEEMsw6D1X1nVQlRiMn6
i3Epz+x+qPmwc8B6GuX/xvInMa+3AXkGnpSyIoakavZjRUlg5zEgSPHxDcT0ryaRAjdrJ9Kwkk8m
ugHVLk/Ob2AJqZZmZ3VwvB9h215T3H2Uxbx5HKeewZ1b8Jz8KyVy6nQ87P+uzt7Pf9JFMIwes72g
JBDVZMAr6658w1NcYNXTqce6Aiy5GYS4xISa6jjIym0+vk9LaTMvnQxKrHhMPhIUMaNd8FEpveBs
W9DNeSghKBKmKS3saPExf1BB6eJ0qiZv8+7ZHi+Plhw2d8MAUdxc6im9td/rSekMAVzqDJILlnvu
GFBIeJqOjeHbZ9XWFRBNQXqpA7J1shVrcnUXKwHd9+6f4UCYGTqPUSqnvKhB00MT+3mSShEX6DIo
P7fGFtLcisEIUGo/aHxtCHmV+DMTtOdxJdinpgvvkBilt2chq+HS3jz2+cO58D4U3iB93qHqyKmo
Byymm5M471YmABWMKflG59r3ahQNc8rnBfJ3jafwdUcva3WS9FGQ3f7m/n26wqvbHp5PX+mKwx3o
dicY0prOkhD8Xw9nu2nOpskdHXIQ39nZHW/fRXouLr7mTDmT5FrfstbckMS086BEp8WbCltSXAL4
aMQxNlJaPT5ccTpUfi8QuMIxNIolCsh4aLISEtDmimktSLXBxQzWAr0FYsZAB1k99KKWRYW8SA6B
tVTB463+Ob2AKzDoDcrpgiYc0YZK2hTpUJ4o/ECDjGLJkU58nYTcSyNcfYPuPrCBR3Ma1LWt1+jE
K20bbfURCMcvh2Wspmia0ZNJ2zvPaIbJLqWqUzcSAcwk7ug2yLwoxfHK5RciEsmoZG5qiTNzXIqk
XYKPnk5eYqa2NVi10Yuld7nDOheKXzsHpJ74O89NyR0qgaNRrTqOv1kDQs3YhVRcw+JK3K3XvjvZ
8tAjS7UJ5Ir920mr2oTtYtT8YwpwaT1FAMpcwqUnul8JLyUGv0LNl81QWGs3enmGqwW8iQtC5qOr
QoIpqPlehRBJg6b9W+PGcfuq83N2xzz6gTwGqcg3HgtZswtkOrjvT0imxIyRW3VU2Om34nlewTvQ
FIfS5hfJfpyeBpYMeO+gxXd1fabdk9yC4Q3t8RptfiW0dWLU/mZWQAI/6ppf17tQLMLU0OOB1pfY
CyqnGarHiCw5Kpiw+rAIGLmiS1Zm9ked9rbSdUfDngu2yngQBr8L8kC+GEUd5TL36FEUx0ox1VkP
L1rbmT1g0EKfTLG6Tw9K+HdxDjleNednQKoVcqACpkG6b2csu5qadrQnhFmw66YTkbfkIi4X5Vdf
BK6AhFHIp9CYl/nA2US5idbrj4WHKa4ahXXXUKQ7jn5h35uEeRWHnseTB5rhDHf6ykqzGKg3ujhe
O2EOWPBCZlHR9uHJtNubJe8d4sDd08HND+REH2ZthAE9X3jgF25e3uzpTBNMWc2Zr95yoK2YK5ot
yCbV7YPitRG8hD0a5eNvi92U2aZBeDtfmmPteyORkiTvMl2ttCFshm3pRvDrnyhH75F1WuImvP8C
jn9zwu/Z1arVj7vAdwEcW6ZDg9emWmsqcY0A5LpBI3UrA3l70RvvKAA+lQVb2VAGOQT6+TBEQP9i
cxIVxzjc8yM8KNqu9cnphGC+KHi9O2r9f3w5CRHKKk09wu5ZZokFwx/z9X4Qu9eKf/p0yyGkIts7
5/X0v22O6YqJgqx3Q/CNkXziRDxvBddIEsw91RRyV1rVZDewGv9zWTgJdAXsbydim5SArkZTQdRr
8GqxorLBl5horUlvR3rsDN1HVDjE6FEmD7mOQGsm0B43NYaDRpr3VkXlChiyFQfmThO0RRjyqqap
9Ac6yyFTlaGIfxQShSRevcdneHkBAYECdglahDI8lAenvQR7H4KDtySaIbDEDjYIvD6PDvO3sC/7
1jMMIV6KmhwgENKZKbkn0gxPPId0cSllpL3nQRiY7K8xv9Zj32mZleyYiG2V8a6cdJjn2SwUWZt0
1VAvtuxIRsYaP7Wl87RtJdd+dom81vc0RsU2snzGFEXqZlHDCmm+RKO1y9pl1fx/eObs/yNvREPg
njJj9evcFHj/iL4D1Z00SO1dI0lSxYWk83A+NsJTu9iZj2GnaWHoBpWnX7iiIj1KhKZyK6BzqOGH
qJIGun9Ffj7+diHPVnx56WxmPQwr7DZU4Q60PaqAfeCu3wsiLtbfTLR2BsTtKuKZ7bXIkBVGAtEV
A/LIK1AcS+9StyqZ44jawOGgmmC+ruVlH0vWNhOy+S0OLPwN/nMxqOP/e7nEQMzOaglRniGpP8gL
i+Oa3NoLaO+rkcda25Qrkvg+d2wCBiYM3++mQjmqPk/aoKeUWoDtpqCFCF17KnLD9tKFCPb0zVbk
hX+kxhpQDu/24RxOirz7uY1c3KG5Zc8THfKmuuTk8UPF44+CnyqoBDyu40OGbrWlCY4mGECqf0Xg
8quvroVltN+8VlkK5hO4xoUygjuXeWmkMjGSSAXB5JVUpgXOtcEaREU8Ebslgzy3VzwjItZhMnnf
INaR60Xn9mxQr62vPwVM6Zs+/s6a+QSSGf6N55XRRAgKkDsmjLseLJraTtiYnpIJOS4slFpdvDki
GhxyiBgd+t9jkarVw+9s5U5Rjn/ijH0Aa86U6O836d+hIMb6ug+Eop4WhmyAByT3gTM9Olw5QeTT
iz+AlzXAO8Fyht9Zucm7pOSYw1ZDraUpBWXS/u9SNdoAoX+DHfZjxrSJb4AHGxAGabCQD3+gLP+f
XZOkUQjsOohu/25CLoy4GqzWmETHmvFtaU4+CvRI46yGIhlDcQS49+PsM/U8l24eehLV0Ic/KCkL
RxwNH+zit09UzoPhYysTLJh63vtDoPHh34H/mF+Q0BxeAz1CPOCwspkYYfQ2GVgQgWFFCH08NwpP
gzt2qDbmaV39+hXkpo3QFo71xAcfWGCFm9ZXNYRm70UjwWOx0XF/3yZgSBJXMAnq502ZUKmrihqH
jlItRWcz6qVU7dYv3xYQRDMbm4Km6GqgKGN85tJYUubF4TcfEbifG56Ym8TBEv0qUWy6/vDgY+oX
ne0jglw7yIXHHm5uOicZM5iV4zn89SkQFKkfReIFacClmgPdOdax/eEWYWKfQf+/GfEUyxwsvd0k
yRS5A03RIsVcu5NZruPlXzD2fmWVvxf91AfqcHlSp5va93Y3QQb7Ilgzf+hgjo/ozJFZu5GgZMRQ
rcspD4oZ3YKX6B9KH+jrYrXQr53Mpows4Q1O8A1D3UI12PS3h3x48zN7EywSayTuf8hX/qEcQinc
pRZjrzevbe1x263OmKpYv7D1e27ypX9A+5a/J+O3aaVr+G1+l8OoziUU0TqTB7z6xvmsxNybzI0R
fc9zuPFVbLZF33XI6xrJWzao9MghKhseS9NvzILN5ZuiCVY9Jeru+9FI1j40hRMyrdpjlmY2Bvm4
gvFp1+BDZN4qORQCdKfa6/Qs6mLUKSpti2rtAnoLmz1Sh1wBVO+z29MOys9f3oa7aWp/s64I8e08
EyjtuSLPbXnfprbFsrB48dZ8ALvFa8FEGzjDOrIzIzZw4sAbbt8Vo9c8HRiaxytC1fL+2WH3dkHp
OaSScvESk+m2jMAtDidw5XKGmtHp2OGrHzamO3s+31XSzQXfLzTAe/wvK4hQ+WNF07SHsDD3iVP7
F++hcny0xx0D0jxx3YA+PnCA2CbRIWiPqF7S3E602WQt785YnRVwMzIlo6vfv5YhGXxNQ+SVJ2zV
4ua0VZ7iJduN9wqEEy+FSmQSyea5lLw/xDXf88UUYuKVRuA/rT2ehWL9lBdDDYr4q9uuLPrdlN4X
f5S6BwCrumWKOOMXDgv+f18fsvf+1ffSO7eLWbLMXQpQOY4Mm8PVavUY8Eu7vM7yVVSIqmJh7Nwj
V0sD+ZH6TJIZk6NJxvu99AHYod6unH1gVhiqjzxuEFLwBoUdNdDoyoFE2WyfvbIofBshqDD50WEW
lVYRuDRw5Y66KpJjfSMxBodpGl0tudQYspuME50+ScDcRk4MjEil+RZzLfiErl4qTjLWTL38T+yH
+yaKEzoKNeupMPrDbX4MaWRn/fikhTEoU4L2JWAgUEFXPbWAbk7y1FA1EKy2NqvlQMaolW1v8ihs
Z3e6qHHADHCa5WOhLSCn24V/AdsVqQir9/T1lRTNkeYx7eQcrBZ/vBTH6n/FBOZNNWty0qMphevN
Af1v1gUMQ0isljJIUlSK9/A//XdWJ1gafXMDeG4bsF8btq7FkGpeerDqoCIvuFpVUmuF+sH4V3eO
/lrzSTkw2xRR911lqi21x3djw8qP3zAMAO9OCbPVNC05YuJrdjWw3+D0eAETkJRVr5x1UL2y0HNU
3zpR9r2IKkGYGjV688xDUChMwDQ99cW8prfNrCVtY9e1WmWL912syU9xFXNtjOq9gBqDG0QAuVIn
Pw5RevojSQLggYS0EAlKrnYb9tp75awGnICc6sknrvFON9vQlKeELR9JgmzRkJrOGR/pUveUulme
mhnZEHlOqeOT8qk1k2lq6SlDcSz1j2EG8wmzGezyc2/ukffLGbFqHpSCrQ1AsTjkqBGeqHCEWEHc
+DOCsJGQ1N5z7s2ycwXSRHjaAvu8QBgk3TvkkNrQEccmNMPrfD4efKK0T31JaJ4gAk4LeErsA+U+
MITXSng9fjDKZdIpfiQuebBsPAY4UzQAwMEd8by9/fu92dAOldKJA6b9hXKqj+EGzIqi9Ej32XMq
X7naFwkDsoFxPX2wpQvUbJJvyAf4H7SN9snVwWPi6xMyKGuodIlDgTchukDWjr0WMDGIlzV4krN2
QcbDAV8nx+Ux6Bi4Gm25gY0XYgB3c7dPWSbqBGCSaYZXqnR5j3sUkKO/bmMj9aCTWsQoHpfzdqjx
/vLYMSENr35AslbiHATDFN3kU6pYgIXRLYIdxGeSTHf/lN/xitE1tCRFk09lLhw/Aj7B3KykzdHn
LbQxbWXs2WeXkvlgrt4qnJsUnLaZysxX7oPxskhTKRc9A4WG4weFtXGHF/bqzP3ojRT6qSf4SBxj
wbMOrJMhLgNDjL+xw7HCIakEmseEvcj9cDFBWMMM3GFgXVhwsFFdk0nXo8l/75Node4WTcwacIX4
zUc1S7D32Qv3N3MmnVWJCBjSEpdCGbpQ/w2Mx+DBSw3Bt7a7k8FNSAq7d7IZmatjSg/laiF3cRbn
wxv24HPLobRIknp84fXJ4Ayq55BQPOK9/HHcVWsWBp2VngUFhFgr9/9ccihjbvKBiHuDbKJMDMI8
7v0j+5v6yFwoTj6LJfh5VT7LXjRu6gmI8azaC4lulfTV6o93+Rmro3G0uXwrRV6FgvxwRNrSo+Vh
D6psWRZPWiKTAYZe/GgOMblJjo+OXfb+he3YydUislHAHzST+wDvcngu7pocr6T1czM7rlO6ai/F
THQIXjnu2ofski8yiq+KzNaSe+RL3u2ro7jz+K0Onq914VI75Lzc7A/6KIegDuzS5uY89EfyutBH
Jo+JOI4i+4xZ9mUT/RZZwqssxZHEWDlI6tnizupt4cQDmH3e9bVlY81uujRF/qZnAN7/TKqAITHX
zuI0ZLg+jYr+M1JwUWi6jN1RgiwO1woIKRKcir29yEog8i0Y/U9MFwRPT0No1/TRet3EveBd9fDF
meilxvUeYQqp5ArD9hpqyc9He4s4nwAq2qjg+tREBwyuQFlHelLARHmUa+riquVxUAHQ1xrJw1qv
xeeJz8dD62XnBHbpZaMtFww0tbn5lruR761wnaVNM5sVNoSgxaVtXxJYHfPdxYD34k/ehuACoJHC
HsoYuXox42D6api+Z/gYLdflBMmBR28ulY7zpZrFv496kqbyXKdKsFy5skEntmOLwwzXCPbW/qqJ
8bu73oJGrCT8nBBzIPCCStcTrRg2JC1HcPKxdfnZhly9vQc036+1B4VKDpPCbkbpOffCmmcEv6Ca
TXu/M/9x28liREeI7n2FYOfA65U33EYqWT12xvLlYu19f5CtG4T2Sk65bHIaOXMTsXcEmhv/wpsU
u1KN6KgCYZruZk1U2d7mJGSamgSjz0Pmb4RwBm3y9b76lko7UxwRUvwAIPOu/6ji4WudAvUGcUoD
Avq9Ogl2HXQSK+hqMpKqGlIRcJayhK9ad+rsFk4SJ44mxY19RJw2kKNhbfY71yUtdwigJ59Cximq
p2A5Wt21LP3iVT213LzZ+UH9jpZKtzzcz9YBsy42UGNfOhxfqnjDeQc2tkaBe7f5+jvCJSKMvUhO
apbyEv4T3hTCtHX7NMTpnktCvBe91KOiDfTV2Mb7Y8fLT1f/gk/6qP3aFMVRQVC9Vpb0ludac8TS
R/ScypyIxAv65dHfeR1M/Eg4um9qW1EdydcO6lKnM8fGkqd8kNadW7HIGt3wMg7W/t6Sba86zPDe
W+/ID5w/pm2rVT2cjHXoTbGcx2EdbQ0AKz8kXupRAOI6nQWB0QtLxHdW61tlXTTmL7JNYijX0P9+
r8/U52TCd/bKNA21UMxZSyZHqVLVSBK6SmCy677Q/P4T+lD2bGCvCdYIpdc7p/RgfoN4TRXUiB+A
bpRxzRMHbw7v0caLUIPkH/BPUnD8dDotue4bPrmOF2ddiYajnwkNDAVijD3pIoS3onGpUnJO3U7g
qAWeUzbreXwkSoJQPBxbgd5ZXthOW6Mn9jTTqFCBJY2JTM/9lVfglvz6qbM/C5QwHJHIT+Hv6Y5p
+4TjJPf4LFiNg3lUootPFpK4+vlgpA+J3ofawv7Xe8aw6QCAHp1quDv60VYVeJUvBj1Vn4FgYKW3
v5OFy46CLdkTZXJROve60OwC7aWbiPfQ7Wn+SfiSxLv+JU4TtxvspBlGCgox/0bAmeuylffZj4Jf
tklCPb9Fe/LXUsxk3FoV5LyFNWn/gbg25kjHuUeZS6+oyAVWfqhUuE+eguxEXCdpHh3afOJG9WLC
4bCTfjzhl3wt0ur9rFtgoAuvK/fhBOtm1NAVoQv0uUEwFoyS+Y+kpeMSb+6IsSvBs4FmE5c/1xxV
ZnUEHus8WwtqVlpGGYEhxxiwDQMyadpEwmahxJAnlRsLjGrHgkcZNVgFx3E09aHNa91KQJ/V49gw
+qnb9lDm54n8II2HWWJkcnZVxnFxmWkytm+Ep8tg4EvIYnk7uLGve7kT3/mJjYNRnfXjlrQzLzUD
8xLH9R0Rm9r+9OPcb8ZwEXc/zmy+DN6gKProkTbakF3f3fGJh5j7AZ6ixRBrOUi46XUaPWmB6582
lI6oN8nniH/uDRvSZFriwrbHJF5MZb0UaOggfOrstvhwFLHGz+oCofE4PkecvdkdzYJ1ZbthNH0n
Zg+9Ak+yp/KAYg4+lNvZ5UDgvuXBBuXSEDLuQIi92WNIu9NqP8hYkgUUXzk4IGJo8gWeaBMISn1e
HvS7SoTwm96/pQkVvdpauV0/R/qFxmH2Mgb1xm8uIiusqIN2RLz6K1Sk6NdGjW1hvL0XZ6XeJKJq
7AHI7WA+Q7rg64HbgEdTh1BQwiY2H/X0D9IpOGXBfuTfE79Nu6EfkApaRzqiWQEbrqt2hmMi+jUN
VWFVHdW9vUw6hQsLiOqF8ZT4d44z57QB6UO8/UoZC21QFxy7PLN8CStMVd/JH5pxaObZ79218sKB
tAMUGPQYb3xyR99gVoD8Vlv2J3WamEOp9/dRhvJNjdwVgvCu47bc0iAxJoMWwCyhC6PMUtizH9s5
4QmnhGA0RlcWXBdyaQHdsbk8t3F959KF2qseahkLlCMfRX+2sh91QB0CKx5XPYiG1CS0EJ4gz4jo
NSzUXAtlj4qLomfxOFQesiX1XyOpjyACZ/pgW5yoFWixi89Em+1MgTURTVKbGR6ELFHCWoqMiqFf
5PNCF7BrNKgzaoUiVG6u8dK8GLvUQqkjA3gSub86u6ZrUI6fD6Y9YfvR7Iy7XX20AwRunOZ69Stf
m6KWEIILenUU6n+/4YE2fzyx2gbFf9dPM12SB3oZcT3b1UKISLyShwho88XRBryxd+iMpyZUnkaO
+DkmXGs3hZZwohoUtICAJ0OQPORrdudganaGCt0hkCwJp6AwiUdLtfSG7Bfr4QtO741VBZUa67/E
/ut7Px5iVEqFCUD3h5Cljm2yOS0e40957UbgdjaZVtDFB5C7+/qgCXyaOvXLIQrczqwTiz5oa9j/
F25moSMW3vs0k3JAF4T2mQDiBp7UYJIDoo/0f9V1zHisXUbOllx3PunHOxbKAVS9E2XxPIc2OKn3
cehsvEfdVHh+5dZokIoTXK6HtMGCIZITVR2kQsTJbyXBHwCekPcfeCoCSfdZhlX/Jhu09Gr1//qx
v47QUnimPkMLxk+6PRHqSJY+6AHsPd+5TyqGDk30amwBPncrmihmqHar4hjpUAyTCHU+dDPXwnRX
xY6Qn120XAFAeTfsCFZrBjCWGnCSCUFWJeMxQzhh92ntH9hdNS94bnXqxemAd9zbmXVMEX7Bed6B
AiK3OOhhVzDcP8RaucFL8yWZBLUfGpiQ+mbJ4uT7oRGuMiWO4AWahNeJudr+dcDOODAuZ0dMnokN
4g+Mf/Bt7ePnnVtTLD7OEV+Dwojae5jbokUDx0sLZOQ97iks85hXM10mQtoadYB8YxRDE1UZga5X
smxJvEcSXG+tufXFmS2UqGkXN4KOb1j8qpwBsTe43OqMzBv8LLX2iDiVJlnfF+RGw2kIhq6leKdo
B4EBnvzxUI+ihpfzaXB4RAir6oaWZn4oI7Hug0R8gg1l2SF2GHXVITF3hpBW14DH3KrbbGp47M26
DFYRd654X54cHMiNkXsuuvAL2C3mtDKXBCxhh6AARNqph9KI9ia69Z8TsBnGX2izGO5zKY79xQ8d
s6Qon1SYplTxKftIz/NhDVTXx944v6eBKpPBjG0U1fBZYzUPA3z8UcaxtkTnZhJ7lOLe8V7JGqSl
AHa13fxA1XS77w/wRNX1ll801CwYPU9RmPzsJk03jaBh4qJmwZU2eNCKLXvfWI2mCwWwdTsYpCRK
mA9b1Ivo/5OdHqc4rklGJmD4lJ41XXAAEB1JMwsZ4Rl0wu3jtYJvjc4SE+NVSs4n7puGadCsODlg
eIPnvSFmdfeQjDydoWkWl5nKcClD2T+De8W1MsKNTNu7AZuFSwqG5qjQDxKF8rUQiN4KlOMKlSWi
tWivDoNeIrToMGeV0sJa7YleKljDwDdhhF2JrJAWDYEWRuMG2ANayD0xL+UOCAUtVrijcJQvce7w
MW43twWzDv7aT9wiIum50Ct7zPViGXwimA4M+uaIZb2lSZQWj/nBuaCyMvJq+X9aGOR8us8DyQOQ
YVA0lDlBkW40ShBOaSda/7r84gFBrYRR1SGm7g8B3HBp+nc68LOFCa0Hp1/TpvqN9w2Q9fqaipYx
l4Hpl5HKLNs7hH1Wcl/cSargVF/cdPmqhNtrQETO0pR4IfSatooqA0Zr1EnQavubxAPGRUKGj+Sf
T9t5JBrSxIQ6RYQH8ra3CAXXZz/0vQ3IMoz4Pp1FRGfBfdCIamxFQ9WkO0hPqaerWKD1a0ynrFR9
sWyql3X2kT9t7YyobTX0kOn4qTnR1oAJtn/sFe6QIuawwmfbzKpvS+uV3VcM4m44ILv7nhjDoZjU
C3t2yLkD6ECR/3ws2z6Jvselyg61ER8meC+wFXdic5G4evroeq39AbmCB2IcH2J7TdfgbZheQoky
lOwXgrcOx4ul3W52V1NIkCCfJy79Slzl7ZNpUJdmDlH+pPpfwvXMk9GgBmK6ToK6EEfulAN6LypY
MTcdYdsG1nl4yyq7hPGZUmJ+VRAhHV9DquaZC387WSuHEL8Ft1aTMr3DfYyWu7mbJEHi2rSOd3KH
DoZ7RUS97nBbdUyeNY4zl6RSzufD7e4bMJ3ZFnbcz6HS0RfvOMxzDAVhv6AsUpUKZ8l4um7yczEi
kXHz4MjmvTZqlCR4Yd4/bkjvj4LSp2D8/CYOUM7/upY3iafJeBooy/UU3+hB83mw+VOJ6i6mE38J
uEt1bBxv47ArSQJ93je4lH8eWKQOvvOdeHz4Rg01MgyV7Fs3cQYg0CVsmt5hEFb9MIzQC7tX2w8m
gA+qIC7K2VOmOcoLQzCG/ThFPwsAc+TTInRrtvEe5JwsBCcgFqefLpRb0IkQQMpLlon+32JM2JHX
P5gchr0sF+JvpUBLdApuD2EyKDYErcffnru7gF6JiR+QaTJ1s0Mp9A21ZpMCZHeU7DI7QcS3LhO1
W2+FLIPAXdtvS3hpAq6hzOJ1Xgv1yWKg753iYxwrD3tq33Wt7pcKK7fzmi6pdIK9TMVK18ogif0A
Xmq7Egba+V5FIXxSfsPSDEnUx70nbmIFXcEkMzhrHOGOFeMdpleHrlUQ2U6KhpZ3BG9qaqeQM+MX
noqaBap6AAFqmrLgYldTs7t69lq8KSt7ALLhQfIqKk4UYsvQVQHhZuogCkER6PleqeKbFLHvlaVb
5Y8Q1lPdNn8vs/7hQMdO00Xfxjo3XK77gPNh6hAqxikjWCUw7juemAcSliIll1i0GNQ71U0b7NR1
Of7v/n04lLxol2+PDF3HSwbJwBbaGSEN31jzRCqn6J+YqK4ZteXztRDOg2BENiHcl3CfZ5X4xafx
Dr9dT+x5naj5VVDhC9/9t52urIlaPurcfqfUPZQXwevz4+QBIjWctzWQ/308SksKDd9PU1l4FGxl
qtagLGC+7K3nUwAhWUw+w4aLZHzL0Rk4IN5jKTCH4MbTQqCuQdleRj0Sm814SHDP22ONJGP0+RUL
JbYOT8kPxwJdvuEuDlJXsktHrT4AHEFDhjObt3DDCO2+jdLWDHyct8hgRNuWeEM4UM6FRj91mDp6
IpLL5JSShAaKlrP2aOdFaOjPPuR0CNw7qTbAoo/WOodd9XUymyjGTUQO2/kxpiiWcAG+pTJcMkxU
fiqz2NcWlWbRT3nt4q6ZbQCke5ruseCaVnSKQDRd+6reTwMwT4BOACnBEOMD6iUaYhVwrmELKB5Y
PGb9yIAFIf2DcQdWrWYFPolixL4RcVEIMzXWrowJlHiJxnhQm3Crikh7oVlICSGsEbDTO8i4GiOB
ygd1jx5Ul4ZQeXtMP+AqZvWoo7PPXdWTHQ35ElFe/kaR4iJvfnrdJs6b6r3X4KKB8m6mUW8syuqP
Rv+FL/pjGeA60yYZ3b9CDpQE/O36CyIBoj9jgnOGZwyjoswXyzFWO/P6dno8UDjx1aoKYO7bP+gP
7jERGVzY18OuNrf5/TXaq+iAyTfh7qNSDzqVE4DpYOhsVkYiA64GbGz2uAciOg0NpMvFWl6pjqbu
Egh9WzoiJnMOWNWwNs2hV6YqXzgnV4ENOimzufkjm1rhQOkrcpG1XfFgQk0CSU3KhtkmXoRxm3F8
yNm/AsLwAjqfHmZXteJFFTY5UqF1H0hzW9KV9241GMsTg+iUtsaUBQGxXxgopIFks4OFrAptoBQx
nYsulZxpYyI24VbRnkRm4dxHZwNp137OqB+oietm4SALlza49HiK2ZFD+Z1t+slJHji4KzlmXM1A
lnZm82+7R0ZSZSAjPUdNrsAuZv6zo4P/b0r4xmpzQ1OEPET1zDGjU3ZOsbDqYt1m8yx6gaay2oeC
ztvoaU8OJhwzhmykW8Sfewvb9mMENxlvDexyWjjARUALhOilrO2yHxMX3jvZkUgL2gtbiU1dZwKG
3tnqmo9UtUqweBBpjQCnsrjtYIb7TpBChPac0YBifeELDic79oeTutrsD92JFlNgkd/SsroBevDz
D0Rxzi8f7PrQf26UcW3BlJTnF8aPvh4N1xB48NvSQytvY6kO6GOuNiLVh41W9vwIpyqT/HMc2MSV
zF3cEa46I4TvWJFD1J1s4itNPvsIpPFfv27pvU/AkzcXRJ4EG7BE40wOZ+v+S9Hd8DkvEbkbg6G4
1uoGjWPtdhU8Ucuow+XtEIHaRE+kBj++/jBJpFUmKiC7yDgrhxJ8nuf6iKfjlm1Jz3Dk3ItY9gXq
sadbqo55Fbh2cHBfCA6QGw1j2nAACDnWMfxcGUS5wmNRLtL66SGHfxIEKNbc/XHGFgiuE+ye5jWm
2ayhwrFbpWMtBTqYFFR3EzsLCF+eL055lk29fxMI3pGdxxRv0LI3R+R/zcwNzm4q+jAJL6VtXEN3
08wWOquphvEuRDsKvnWZcMhhYw5HBW3NeoUBgdlHzV8PNYVqIuzRRwHiVocM+Fk9vrdgFJwGDLCn
Idswk1yb7aH1folS0Hm3XhLtbS1dO3bI4ywRqqt6kxgalQpQuJXcujVkbsi22fgKadg6J0P4ubmZ
5LeqP1wfGsALKBKTOz7Qs9zW8fcnuJIZReHfKG6Sm6WBZj+xHXzzzX8Ssq98+TkrUQL4DaUG5gFU
TqLpxcw8EJFbVC79E+w7OpDEGnatW2AsI7xRAqNOydIUqFAjzCOc3gY8rbgChIPA+OM+i0X+8kJl
ni+Aice2ZnDXy334M/B6H9oWqRp4NJJiK3TqOALOqi2vZ4QPzmnOk1Pa9QbTyM0xB9R8n7kWgA4g
ofhiN4jlmeckdhZRG+294qCLp8caKES4acrLXacedGJz7AqrHG/OiM3ZnWWLx2mD5eOIMNVFOXQ9
rY7VsBCzUTxFK0sPhroTDx0y8N2tMMxHA5VR8C4PRg9ziyYXWyxd8+gAU6ZUJwfiXPwnKCQzYzic
N2cqZ4UvbrMpzLwsEnIJ85+9RwQrrVEz75XjiJgWMxxtZAhoYnw2865b6mvUVT6BcC+M19skxLQD
05zvCvKi3cZF6Vq7Zwl9YCsNYTwqWb/gVAnU6Yf46KipXtRRGCjuHQa+ZWbQN+7XSwllYmqyAMGv
d/or1LsmEdE+y8uPcZp5FqfGVwGaqtD+nLVom+aGG2+fXWmKyvQu0n/C+SfeNj+qKVPCQhY0CRPf
7qRbYRq/Ifx6+gvdA3HwxMTQHLptway7Zv38hfVywcRmX+qyhcW11I+oQN3grcpxL8OQUov5UDov
/mr/mz6J93r4V6/aIFRbU4eQqoJkKzTEx2MFfQrDD7aaCxNygWVrTGlp/W5Q7v/aNPqEUPoqxNCl
D5xAwKPHmaOn8WOYM3HoUh/HiVjLg3jtSINCHHOssZBizHl/FL87ssV6CUmpozEnkgks+FUka9I/
ks1AqwssxkepLhYk9wNEPSfA9bhsoabpvDkni4BCF77DCHNzNPxNdSvgC65txqYCc2YQeOrKI78l
MLQmKK1Bd2hetY7LbHZ8TniuDmE7szJOfCanlttBsYSGzqqQV4L5sDugy/YBkjumumFunQCiEyku
9U3iTsoLRqqisLS6ccmX0hEB9DHf8/KOMSxHx9bG+4/y0IDn3yUzIG8DJhnSJQhmRhW+MMNqHim2
C39WWHmDMBwldhGIrIxk97oeOuLDq+csdFjV1ad7KN7KizC0xDtj9ww75scvBAKJEPkgUohvOQnj
3lbeLwt4439ltPSDWFHu+aZ7v5hCY1L7WeVj5aFG/jfRylh+1VLO2pq4C1ADzhG5SEJvvmnXu7zK
3AALkAQPY28ktUq2JxTOjxf6Lt52shfs3MMDoQ0PHw0h0NGoNZ2+RONAYa+RDO7k1sRF/Fso4tky
kIWOOcqyeHQ4nYIkM/cBYtuZhTrfP9RoSiwEESnbIGOotEiM45EyO/l/tY89hBL1SGJi1IPtYjAz
Njjp+zccdILFxLAxqnGcbLV6ViciHu0GnF3/G0i0NTfZXW3xQdj8hGH6Nvw2MjUDelM78/+UPrSU
3blvbX7dV9mCyXT9Z2HfNDIZWfDNpZEcNngTsf5G2Z9FXg9Hppm1P8d2tBbLsoeQlVX//pdM3UZn
XFEObOD7yUTeWsLT0XwKFdDZkSds6/0gVVJv5tSYVM5gUBPze1qsD+vG+z4+A9Z4ukA2EkPtPLfA
iiOZK6ejIOAToCwGibAlGxzT5a9fSyRDxgPCCQl91oPu5vO34vKPe+e8BD7rP5Oin4hGhvag+sb2
b5NyUA6MWBenWpU/0WW0Lq5xb8sP53kA5hlBuh00VTqp3W9PzslMgkigi43mnOOQcAPyr8wV4N0U
WjqfOqGFKaHPeyZ01sQtX6wVQRPtv+JeTftddZ1bndGbEkC6TEqbh/llHy+k+40S8xwh5OCYY7u2
0ACOSAYsGLgSSdOXdryHmXiWkazkSSoyQfJ4LY+5oTsjKjFnSWfmYBKL78ICc+ry3TqfMbGr/E1r
SV5o5lJuh1F4FeEl/oMXPn+yvpmafgHgIrDWW+XtXOGogh7su2bCIko9GBrcGj/fsarY0doRBMiu
gd0XKGg/KJMolEgyH4N7bbCC2PsDOtHoBxsI3hG85FMv3ci5/Yml8PlEcc6bPEmi6S35Anosvgtt
b2wGE+w0/FDYKYGtdHABTZXWA4QZgr8K+trO37Sih2nuIVv/YiebjDRumk0qFn+iYEuD9zQVp1P5
KVUykSW9KzgDf73eaNfqoZUxrWI6uN+5XEKJzKedZ0JFC3zjQm92/pqpMKIARSGTAh84N85fb/xg
W5yJFiPJno9woYF+QBVcSm93RbrVkxVjKZdLqCTUuofcWwO6zWe6wocT7ibTK7CC+nV+7AwTsOov
otEAWqR2r6Q+Ibm2svL6nKV0jbSmbI+wf3nEtcLkjB1KI6yLcWO9EiNWb5cqKqD8hmyqF2s04MqR
QywPASy7W0QL/NyHuxe+NQmIfuMfsR33Z2IeAYDaWmqsQ+Fh+kOEF/OLA5IBZrzTL8kkso4Fei4P
wkkKdIx3Jtt9YD5HFa+QJJuoe/OVlEZM6I//cUlx3B77tXT30rIzmIDahl6Mmsic53Dne+DIUgtZ
/8aF+R+iwvmxlRfmNnTVN8R0at0aGQ5uTV4nT7yv/9TY280EoI16EsedruQ8ciSxsG67ouvDW8+2
ZQZ9dORsXhQw2zq9PUuPMJMuN9vp8Vfr64ZN+fprbPGSvN2ZsvypSc++6t8Qr/mU7WoVgMPbnXxl
0xg7+A0YgYyj2/t859/9qIylM4LEpOVltmTQiK7VwDcYsoW0d+Y1m0sSnl5BbZv/3GgvyPcgyzS5
6GbzKS+khF86tTl7TMpFU2tj/3e34CnWLdTXs2UA8cpa8jtZMmO8vyeEQcSg6sJFZuDxydFv1c0k
XYJWnIzMBlmVDnkr872fPk0FD4VgIuzWGQ+GxgmBtlTS6o9eeWBXTknh/+vKVzvnae/lTp/VAoBV
+4bexZjd86JwoDLm1Htb/XockJO9SS6p5Z4pbokAgYIl+p21Pf0U16BtkEW3bqg8j7bIkmumcWqL
1ONDyDv0zz+8/E14Wg3QJerUcaUz3pHIJyAhEg6LBQs7oMbF8zWMmYQVyZdP/bk4kIIclvsn6Jlr
V1Kg+u7MQwjbiq6nu8QMF9JI0zytU6y/4xN3th5Luf69RFdx5kBMhMh7EcCbJC/HaLpOVMIPmsq6
Py2XcYQL6kiAimADVxzZYJm/vHkjeKuwPdz/6rdgq5nwnSSGOCR3L7yeBMZwLRUNpej7TnzBkD61
h4q81G4q4Xw1MTfBoJOVaO5ImxMR9qmDsxQ5l2jIqEykwM2nL4kNWwPg2Mjv+XYOfG3mnZh99Ohy
WoVHw+3VsFXOtNHhutEhUOckI/72HajDX4fuw6/XKh9PAK56Sc6KVGwvKLkYHL2loi9BaUSE8LGJ
DNRk8MARxghmdgMD+4l76WmAMIcL3qq0JN/nbBvYYC7AadVwpjzHOiGgVVCZOBA3Y1E4+NMa7VY9
CO75kEPtZdX8Qrt5FU9t+9BatgHTWjNt648ny3weK67E/QZBF0piLj/hFvuY7PfNUPGOTgeMQy6O
enOK2xssv2bq5iGPjXwwlQ+cKwfuEU/CAVkJlDfoaF3I29zRm2NJJKB3hN9B0k90hmclMJp6LEBu
lO6bqbhuLg/maWD7QcUz+SgJvWZyHUpDZLMR9wVBfscdX7GH3sbEZOe4Sb1MqDnFbm7Ty9u1XX7v
ynOxJVvvi4i4rDH+VzKWIaiNPXU2HNyBH7bicSzDkASVeR/AQZtqToc3tSIUkr3jp1wN4f3x5gu5
a6QgX8/yns27ECHvK8+CVg6CT9pZ/hrwevwcEFUx73WMmd6MHlXJifZlosPdTIvY2IEhS9SuiSyb
DNuffURcmMp/fnOZzMc3Lc7oiRB3eWN7ERRhKykWndBfRlr+6X3Ns5biTlLT2OA2eh5wwV28eHet
tTF6onLlQRfnQ5eWu/aFwFj+X1huqZHAMQOSaU2aYu3LFvenLlGRKErnB/pWgQIzILMPhEQEYoNK
TnL86g6PXCkpQBeBIcCC9cg6VQ9GqpmRYRh5Ion6d1a18UwIXXOHi/3Is8WsX0qgsPHPRiNRfU9d
TvGDUpfHCpu/ANzWIEaJ+tgWOhB6JWg9GSFnSYrKJJ1Llxj/YAaChdIa16gR0Nfh+2Z6eZ4Zsqu9
/QOCooNi1e7Ml5bbWKoz7vcHptzzwZesArP45GtPM8/s3pUQxagwX3K4Q60LVz2+V0wYPvt828ur
YId2Snxh464Y0+VCQRbDG2kj3kF/Td2gxqLVUI4HBi9/7yzlA1RB5V5h2WhBE7Wl0SuSprrFouRE
EIMBeaYlpXolxAtuGUKtfTCk/K5X2tHdhT0C6TUa3kQTEJHyGXutbnMptIqq9GCNnw2lpmtgoE8w
EhXxj7J21DU66gy01OFDwdznw6r8yfDnwqsUzjEcUcxHUMaeP4nnuvZZmxobFnbdVo3p10AoONlZ
AA/Dsp/TwpQhfHVq0cA8vXL8NGAbi4lz/TdWhj7eZIjc5XR/BGzBrpcupokIn483TAlh29KoKFbZ
wV0f8CHc/SEPzIcHNS4rp0HkuZRbM0l7qntPIpPVXwHoB0A46SOhidRLbuul/RuEyGmq3PEdBsNF
TmVjjRdtF7XAq1AyPOG4GlbshJfgbLVshFJwrGNb5xGwZ53r0ZpCG2e23et9Oxjr7QTd/y2i12ur
/kRYkxJ8857Rc5BtEhTtdFk9INvM1SA+cs9RZ/nbXNTHRsFWGkHwrxbcfLuYpW5whBgaG8M3TpMc
yCKxUdmYdF0nR6ivXjZzigfAlVbYjvR7q5wwTw2D2sZJJTrwViScsPYnwBscnbPKFExQnomRDsYe
uV7atb8dONEihLK19w+PtjxUDr/Hhmzl8SsIhf2BNtD3exbTwB5zxUjp4hrIjLC4L88NzEu7NltF
0un5YEbxS8SK8vAQnVwja2rbSYnO7ODSh0x+EK+s2H0qlYxmA0XazlHpiSddtncQD3PsqcV5t8Qv
HHdrnAOcrlbggdZFUfgF/BD/a0v9V6fFRC0aIf+1jQzYanVi7axRw+W8esRwbdXrS7aaxprVFD9T
Xb62eHtkhAQtY8g5ucgX7L+m9rBo/rAfZ/QB/jAW0L0FUu6EKgi3TQxxFt3skcxpkel9wsl3E0sV
LnB8GAb9Fq5BG+8VNvA2iKtRevAVqa0p6cK+vYgtdRuBZZUnjs03f2vNSGW/m9n7N7Y8vl3NFw1e
fMG8iqKWT9boADIvKZ1raCt7uQue1/8BKztq5dtwx8TA9cKZosZ+G7ASETPoY3eyh9TWaQhIoRRu
SRjoWpsTxdPb9vqaUJoFEElVaF5RrTALru2a5d3UAWVCmZKu++Zy9mR9YlUza6Ppy/yLfFFc8jxw
hF7PtrO8TV8g1q9zwrIwF4W28qEYk9CbMNHC9VGSc9FpZnDIruThJKPxg5S4N86ZRhisM9aEbTK/
YsDL9IBJuIaZX3RlOA3bMVmOI+JUi/BlJsPhSrJGUHUpBxz637j7R7sJat8Vq7WlFw0QE0AMbb22
zh1dw92NbnW5kssB8611jAk+UZLdweweR1s6Z3hfo8V5UR+AIFM+BykYbrwX/fNTtraMN7FxK76I
mtRenXq+b35eHWgZm3R7NKYcVVj5kDalClvMk4d972fJ6UlBfbrvehDOqsGT2ONoBvrAjhfkPTHL
0S7UF+vJ9TEZHtd7X0+ZUiDkIakMJsyIlo5Qyk7XMeL05JDcI5sAVJqA1CrzwP70KK52vyrgvEtz
iSoEErG7cPx9wUVzrLmkbqBIpF37Dp0IhcOtr9aO9CZIoyTFsFrBMfF0NsiQTEJR1vGKVr91TKc1
M88E4VUi2tXapzl4eUqSuKos2e2LBnq9bhzmL+wYVDLkL5GvRgRr8CcJ2dm6TQIIxr2BOCNLImhZ
X7ePudKTkvVQnbJ4eZVF2Jhr1Qj3gQ95d8iPYL1A+FO7pkJu0+NG/LLJZ/iRy1RxDYB/o6OFPyc+
pM1faNQyEKqiYeI0pryuemtuMuO7m1+jLD/0NLOxBRcrWjd32zzhAyaPOj2jON7oCIJ1PBIvxH54
HYz5axK0rvc1bby6cqXGaazQ84kgID7nk6BqGsEyArxpPvN5kctvIFlYLzvMZT5x3Teuw545Wk6R
2SpKEaloYnTga9ZNc5Z8m0eQQ9q5PdK9upH1t67VenzUv3eI6xCYNF8Ln/UBZiD2ohshAAoumQcr
n3DxAj/uNFxiQf7JjBGDa6XIhjSh4jwqWJwPHM/FM0JW7X0J4cXMX1Ce2ofdfT60EBMEIVdizvVK
7VHSlR+SfV5S9TpCueyYYQF+Z9Qx6ly2+wYRmC9CRVXpYpBmEmP1kX2xmP/lBhFTlHVb64ud+Ysx
EUy7tZ/QUIb1cIDjm4yL8CzFbPQevIXZE798z11gh3sNDK2VMY/U+EASYAeUaM24udUAIvnWolZz
C6p2yjHzQ6WFAbRjITvL183OCF31+kr/El+RDxTBAdPWAlbcjf6/ex7yaf8wPUZVODnEmtZVL10b
jhjd4bnMR3sqC9Q0L2FkZavTnS0uM4MFmgH5nv6VHeeWoLTOq373BT5s8e/USVucKSEsxV7vFQyJ
zIsHR1hNAmi8m64Yp2cPQVp0qr0m+WAdCyzk866n7wKd6RHpk5cvRZXNTBWvmhWV0Kf2HUI863nY
EJlLws6hdad02ADHiz/F40Jz08IJ1pj3h+QoQ+zHonRS+Y7vUwByPUHVG5kO3BIRBmuAIm/icFvk
L3XYvJEJHnTLbKu6zBM1NyZgmbzV5R93jE5gokGpNj3Wde1HyA2/gJSjHSeONj1UZDxTlrCGQKhU
kT9LtyNdTwMEJXJKQIXNMZbKVC96HuS9uM+QfucvxDzvfEIl6ErxKzZwbPGQCn2FgN6cgU2kQorK
r0pgX0pf/ftYtkQJPoCh2y9VnAzgzZf/vWCXn2wmXTOtK5KYSJPl6ZbxvwqmHQUm5DPbBlzMuhIA
G+KzK3UpggBCkAmVmEEo3P8eVOFBCz+12ccif1ZqB2XAh/+v6UxeLv6iAnmvp32CVNCFAiI0Kjtl
kpVPXTSEr/DUqruniai05I8adqM5ZGH8wVdM/ctDriA3RrMvMJOHG1yW5KaFFRUMD1VYUPuq+nnI
BLV9hf3J/cRmH5ps6Tbf79ffgRg8hskhE8f6BXp0DotuKtLjmT42VA9OkZ1IgxH60cX5peE4B7zz
6O6DvywdDmlPUKrNNPP3CMewm+nmyDFjLtCbo5OTwb7K8d7W1KgCDBSAt9vVZ8IqbGNGWbYl7seR
ZsNtb6qJVD1qq91M2wpNDnCodHHs3RL5J1bNz7cSWkunbSMAaB/GDmxoU2BrmVrBcjBaFtMtbLJ1
xNvpM7/pd+vB56sSYLCiuoIPPNSnPVhxgatjAzXs4Qp8rMYITE0ruWfagjqhBOVSutWxABVVWMzk
Nb0k25LUeQU8gWAMAWKgseU2P9RvhCGHi4YPm6n0DCSlBfVfCEVInDZEVmcLUkNK1n73vX+GePIA
AvxalspvpZmazruZuYqzHq/Z5NBihFoPHnHhXWZ1bzoGytTEAaBy+agtIBJA/9lNXFCeAM3SX9fh
yRJnB2HPMgHKQ/w1AJ3TkmTu+MytS7gs+p5piyL9djm3f0P6A7B528cXMZKqaUgWqxPzrMu8bsv1
dia1AsO6PvYqiwSY+jL1kSXGNH5AKn6Hp4EzeGxQ6lme2jSW7hoRGsVOAxqmkW5iDqvRaxEBciAY
yNlqXskDvoJoFRK9ddHm8ZF2yZ5eLt0xsABJqEx8Ks24HzlooGMK7/CU5wcow6pecQnzVfkkZTSY
A6jwdBhL1bWhkhnjDfww/dkI3u0XbO2qd8RxvxF0bUvXZ1GenDxpFiq6IylT7m+YitpkrtNDWLPA
tWKdlOfHrPlsjCk8z8ev1RvfY6mxy+IGJdmGWJ6aEQYtpUeEBXgfwriHpUUZtG+49KsIaBe5gDDs
4g8h62BbyLXBpipjYQG8pCwvxeTmlvTlq/S5+KGcK+fP4E7BJoewvNUU+EvWr4jIzC4r2BCRm2Es
1SuCeO24v4wvkHe0mz12DDUOPfXTACasYVho+9HX86+c7Y9VqhO12EQ5RQIIPDdJ2nC+qlcrwc+y
vg4MKRngw3OKhBkAkpgFuLLvAk9/3uJ9r38NdzzZ9ZefquxFCPs24c8ohHnS4zoTbWxo2EFjVwt/
qsTgPY5K4ewQpG4O3WBioNo72+C0hzAX5nWnNwCXcdevI/hM1Hrz/5V+l/ZjCz3/dXegpC1Oh4P8
uVQ7CEIGwrzjawtaCMr8BgaGMoLZyBt2ulXiw7g5b3/rD/mkErIn2kh+brjlpt7bmNi8SUoEeW+X
I7T0kZjwDTmV5V9AvtZlU68OpMylR+tSW33rPOMDemNkrfQI9/B7YR54fQzfSO/tDyOAt7uV2A9M
/HyhljDRSj4dw9mzF62KDvKL7bKelRAa9vhisZpnFTSSuNfhxgJb3bUaqDEBbp06XXBHkl+Ng0fl
p8FzoxtSPwm3b6nmg9cz3yzesF9y83Mtl6ulqfu9Sl1ymthOI3P2r4jq2G2UgVm1clWvKOErC2WJ
6yLDJLIzXW+m7q0amjoPG0AqdyRoDIAiZMkAbaJ+xJv+tPjVupK6iU5Zet44QutMHEfSiAmQxlS2
SO6VyUvymnRxixXQiaLPeNzw+eAa68VJjXqlZYrNFW2hYSVc8S3Tw9O73Nq5+vvElfX6nRyMVIjr
crPvVQeB5k3hlEP69XB87MY4oU9rw6h6d6WFBvd1lnZve0v3dkfwT0EuKTEf/gKeJbjGBZiYegIf
2ch5IQ35lsA2WviFyI3Uyh5Q9pQpIilc/Qnpv6MOlWuBmd6s2JuLwAXfpZ1sR28CeBBKoNJiU4Ua
A4Sg+od+s/9mXivCuJL1U3/b51ydj0Ac36VgK3nuHWs/nW3grYnGMyClTXxKyAKNF9WvnaCBFgfq
LGe2bMf46Ay/2qK92qSso87TGLnGLNGu9NZV38+kg8dufvYpfNmIe0aSINrdWdhUEzWrbZf30GQS
FXquVkRowFQIUdx1ZdhoWk9wkqqZED7/YaS2KivT++l/9CemX0Y1TEYwVRVtyELsowl1jJBTtYa8
GtWCVXMNqLHtO+NzyOTZK9ZcjJVvVT7Jbpi1WxC0BSx5SbAymG1b40MDAFyqWPp6/3+LsOvSBEOG
nTfyo+WH7xEhSTvCK/Q3DWehowaLl5qRr+c01QcJ9lOfpzTh8Uy1qXlL3ijkl/AndIDjjNqaoeH3
SJn658cC5sqzPjKLck9geB/N96aoXH9UhjfgB31DZzYP3pQLCIFOkuGb3ClqpSmZPkqIDTXVRIpx
Qde9mXV87CE2UTVwIDNgOLoYYcqdt8xpHn04MhgMczUV23JYFLNDERqSQ5G8td9Te1Ms1RrNam+/
dFEmSTQCe8Hlb4xN+wdV8d0g/8LfPNz9TrjIXZoQTu0MakWcQq9o2saVmzbojY//i4PibyknlE9L
80zVzcHhD3hnBjlW+36rfCMRBdfviVf5BWZOQMmByZPu0ubkHI0YGVhMOjJpXP1wqINuKQLLUft5
W+Q/WnAxlnLkEk65VZnSWF8cHBje+hshlENZGoFLUolCo5Yk/Z6GY2ECZvcTj4WUd6uxnFzEwrft
u7q/Rrvg4pgPvoD/CUSM8idx3TKdLuJkxu2XJM5nImCdVsGOsNRaZ1c9YW186y7hhdAJa2fDQOY/
SbV2PEaL+Jt4+qem8cJQ7++PYWMplwgEBmxgilkwfTbWr6O0vxnncLoqAVGoDRXnWbkjnFL6i2wp
tj1MU01LeoVnazEcZ+Acldt6dt0t3wcIGzJri8geAx7i6/MImu4cYKw4WVaCobmSnquSPBqPd1hM
bHqFv9ITZ4PfjAlNxn1cd19DAPcDKETGBeiEGaxLXsfn1ZMdCwRodse3ZIHKI30j1zcqqGy/gGta
fRCeM/jZ4H/aIo74jHYNJxpMGUqVwH2BSf4ar0UFxJS0b3eH88FCUX6ITgMPDjdcGphYSQ97jdzb
0C2lSiWdqfoIcPpClU5If4IfHDbdiiaK8bF+tz057/VbI4LHTktl9zTrzYSG/1zqdqlOofY3quBG
LDz21u1fTKoYGEotZ1iaAZ6bgkOrf81QXrvt1aAUYpkvsTVas+D1M4tI7i3y/wxEKIX+BH8fH1Df
mlyPsI3Hr259uIX9tzyBExARciMOH8+ee+xDVQky70NzA+cfiEIBP4E2qWueenbdRb1tXztWARMZ
gdBL7SZV1Y+a3n8NfC/PoWwPzXMRz0Dni6DseKluix4pYXxfBgbGDKpMzQ0coiHHUztNYqrsg/G1
VHbSOcZ4hayK2v2UWUHSc0392gQDja1TXdpvebCq5EE/IikV2WBXvJOL5pHaUvgI2AiiBMB0WVTV
9hVuIiBiCohM0X0/62Xtp3L1kIG1RA95pES0JY+7rwQpdvguTtoZd83HDItkZTQubjYiRSEJ5Pou
jBQ5z5yD0+44nahwsSMgjLeyB4QKZSgTfbfFrOz5heEX49dFMgJNmg/Bapc+y5jiA0Lvidi7Fyb5
hDiU39Gvadc8hWu7OW+TzOLzKOTE8/+43HAej6dy+UsuuH+rDf8vm8RpAIwBULjXcxYH9SN6y9Yn
AimI6DvRsTB6RyA7j8awUceHZ+W2VqHLKBXU98OOPgP2hAqyUtvlF/W/cuGLbbE/rdRwFTfS2PUU
AsltMNtBvsrjKHdgZlxfk2pcTj3pXiwwMjjxDwo4oF5dIyURPMRiYWStnzVYtuPXOOCfOlDnPgcB
e8s0ER1+P//gz9S+OIZ7uS8N0UzDvR3QPk6jyFIkBuP/dUBa+wbRC5ybz/clxKkMGDhBt+5N3HxD
Iu1YeIghckrY5djoYrRSWvi2IWhHeNMXTtUJWa9MTi6VJsfznnwvicuJehG0kbQ8iDxeAeritOgu
AkwxqMLOmUSnPOSN+Ee1vQvhU3FtAjDH8qqVXCFABML5ltExouFwem/mcnTz8Ywp4hhayGguViYg
q4n18eGSYTyjaP/DSJMkAQwvCxiDcnAZkLehGW5Sd9KoOd5oNGj+G0NSsmuqp8se1Z6VkfMjRn9S
Fp0AALh7ivOS3Cpc9PyKZ++zDDybO74wVsyZc++BiJyn13zYCGikShTuBXhwpEzL9ocm+gDag/ow
f3axP/5KWGlYPhJWWBrz/AD6JfiYC4ENYmZZ8YaH9UCAxO2qJz0msMqfI6H1KhxPRO3qXmDgM8vy
1uPDnf3cpoz8AqybyULx/21BGvtQ6ODDtdoWxJGdncZzQwLeJrSTV9n33oqhTBNF0R3PHgzL70VO
6a12pKizS6SWXWVIoWf5ZbmhZ7edGbLyCXll1kzlYKOKbV9n/jekD8Na6iXwvc1ZFeF+VIrYNoDd
PoSqjprlQZ0q2gMZykEJeEdWNQxgzmxsMXmV14KolNUd4ilvYcGR6nJCw6SMnmCsiZqWzg0SnOU5
5o3pURXfy6tHPvQ61RcGXWObYOBpmty1iP1JU/rSYPVwaiu1z52oR0ecLfU+zfKRpGKEz4JaLtBU
7x8EiA7NJXBEcqXOyDNhGyopgzPf13rRo5dTVCHP0BRoUsrIeNMAHPRRGMLucMWr1mdqjNMcgBqR
/9atSqoNcqIXcF7qNm4JVjVROOwxbr0fcd4SZoZ4BMdZ0YusMlmkSkOKyOjHhWBR33QvGVUtWQm1
IsaXhZZ+SvjgsYMQalIiL1iR1lXBCVZfI4ks5xhlUSAjVI1CpuJWDqEhJ2+C5QVDXa6O4flP5yAc
AwZI/ivUDoQFUnWi8+kLuw6+Vvv7feC75i76eN3AuJRsuRawbaR/lTi6tZzLR9hbEJ4ivUPn0iZ0
dKJxrNkGgClTimoRnHfWtIURQNF+g9yJIxxTTgx7su2/CmSklO6TpZ3evY1KSwZhXMsQ7/1xebqz
TdNFBaeGLnKMNirGYZhTRGGUorSE24pBmGV0EigDfiBTvGca3S+HEWmcTAOu1Mi8veAJC6s/bgUZ
F8jXZZpbGnbjMkrHzlNLL8KNMajDsVqFHvGpaiM8rJYlFstZk+Rxs8F5yc9oNWMdoHVOIrXvpN9c
hfdrW4jKCGK/m+PYgOegeAFKsvqJIT0/+Lahac3H3VldAzbqPHTCAhXaiuukK4+1ko4NjWo0cq2N
qwA0oAxAXNzX7VmlhMip1ycFnu1XEqnxs8jcicOJZXgNLVlVXnhU07XXM633RJ+jE7YWGmkWB4xj
LUpTTMUNRFeAQd3CBND31R1sAH4SeVVLrBHKOOG2OeS6m2+9GC6598dR51nYkL2nr/oJH/u3cMcU
k2BXIHr+RuXF8wI/vumchhycWBU0M+WS4QN+m6NcK61o+OOHimrVTZMHckFonvvjBG6FmRbdzAoE
30pRwTLQgkkzCnc0K+5SEu7TYckMkJkj6bMLodULaEvlUmr3PxPoEQvZttI3cuWQOBiNdOIX8c2Y
NixxjvPcfihnca6fkqHwPqeednV09iUJaHOGq8AU0h02uC64clvbS5Gm/9VQqdJgkeEz1iv5QAN0
yfH59o5azxOcPoGHyGuY58HcPVXTWF93/N4BBOWy4e9+or6/4COX4WQtKWxsbSDWJ5ll+DQ+ZOeb
VsDbYfTyFOBCRfdAU6GgJka/uWqB6iuDwDYZ3i7laqazhbwqseu66Apk2f7oqwymDH/bGFVisAeb
qmvx6wdwloStliYPfhPW1jFQiMIJy58SQ7zYj/+eycLFhSB4Cr3vTCfJR1csxwCOul5/p1k7r/El
7/In/Y0Nit7BGAaQbGUl5094t/qmdDK11IhQMIMPpd2m5c489VIJ0nmsGzkMZHhRI112yRdiZuwM
LRNzOeFWBcr5kZceBZRAaOIgwpJUuBSZ7Ddmna9thLt1UN2hLpqRN8N1XI5WdezXONUw2E2R28qW
5Oiz6hgBaoKqSTulIix+9+wLQN8txauvA0LFwer/Dl5e7t00o0XgHt6K8jrKngkd3DHKj+uXa6ew
f85qXBnusSVJUqc7BFq41DYycw8dUT5VxONcnB6VLQjl1h2slb18GhAbldNullHiO3K05OX1DIj6
+g3u2mFaPUIfWoDv55DXodcrNd+amrrzUGV7kqihvjM3I2crPzFaMFJw+4CtxroGYNdSoT/UlRqB
mjoJIwU3DPsTI9jiDPejmkgMxwzw4vGh4YfnyvU35XSToXE8biVFewjMs8ftn19DacX9g/ce50Gb
OhljK1BpxI4ak99VmfJhSMCyxhCBcvsBU3glRNSK7kot/oNipWIP1qCVOCtRpxkkYDsCJMnLbjJ9
DZLlwQXkoMvcGZmQUqFgThmN2lXzudQRm02miwZ97W6RlBBlzhD/gHyAxe3Ib8dMKijs3K3d6S3G
+RmueS2qqbQoH7feJxT2jOghNwtqXaJ5aZ/8eh1vo9lP1vWWEaDJXY8VcIxa3bMT3Ifg/HJZxpfy
MeIA+9+RF+uHPuezlEUEs4204DUymhecXORX+SINPWKGE4AgDe9i/Z2VBzEevpfWFZqFXbsWg7vl
KZMWPgeGnuedCmgcHyHq9yKhxYWJXFO+49Svf19J1X2rChRpwX56kXsbn26CVM5xzfMaEQpwwF4R
C06+qZQOsijo02+xYptQigJgNPL6h4QUmsakgLcX0RpX2Rpmwtn/U8cFFP4guTnbduKLacC8q8Mg
h30Qyh3KIJE4PReGkagqL+QD/M+XMLRvM6lfdP8rbi7FY6XQghh9yAGv0oCtPfuLLx8mRnFKyePN
oVKrGeC8hJCsDoSo/rWTLUc1U87rKyNfOL3qSh5XtihIYlWiR3elm9wdbQhqlaEVBW4OjbcGVEEw
/PiJXkD36xAvfjR/9GJ6ewHX2RpQXuER57vDA28focCJp4DgUn/AOcVSrDcYjGCbXPZCY4S84o5E
jizN69q5d7rAdCdlmOSnxbCHjPcFIf5/uIz3lQimOmv2GSoTr8YQTp0s/siGmP1wlNicei3p49Uf
Yu/Wd/ydPs0CsWeahr440WozINPsONeihECUn9D18Thtotm6I/28CO3QWlgZzH+izUKOHbEqSBuG
WWSpkx/ncgDIa1P1y5ZMwZ5oDQPZtlcEqkP5NC1H6jA6zLSCJKawkfGVago/JdlTar+Hy0+Us5fg
7mR9qPeD/XqBZ7a7BWss757+N9UzTZeFcuuB+l6YLtLk7iF/dr8rSNVGAQhgB6gflliwb0VcduCD
rQpeSTCyaJ+xp3qOzQqVoknWgrLNhBqttA0fbWK88OKNcjHlnnyg/FB8L9T7xnbeD6POZltelj6l
zRKT1MP8hPe31fPMzdDEN1nVYRtWLtaH8vIFFQnTkSe5GwtnBHSrCsw+6AW7ysSAUPgDoxpD46VF
sMYGVdM54yHsxMH2igXAEaXuwDoIfsd5+ezrM5sYktbk0RUZyQd4GYDewi7o2LX4oAgTlRrLe0k6
K7AVqo9t+E/Z9ad1o8tSAHZH/sKy1DExMmA+KjxYhoyQYjbrMHzRFH5unN+sg7NPGZENvC9NF+Zc
qWrXD6STvw39dv6vfj+wdc0Yw0ch4g11K5bSywK2vLbwg2WETibyi9C6VharONBuJcgsOArw8kxL
nnyU80A1KFrnFumo13No+KQXEG3YmdOTWr6jqIQNqQMi1ChYxSeXbP2Ex/bB6W7vDWeOD+hP+Zxk
EsRpz/CJcH+eJHgzUrdVlCXJd3HrVS99llOZdnPpFuaZm6cNqRPKhCF0fS+YOYoRRs12lBU1XebZ
nRtu5rmG42/7uPSXb7aUjLlGiRbfmLYISE0shoFhiDQRCNmTFpiiSLpeNQcezkNcFL27oNmqPNZz
+hBr6K4aK6/3vmxgG+LgeMbVERtMqLcN/sE7qVsxlCnbbyX4yBTqvOz2wp+Ygoqm8/HUbmgVqdNP
9SOz2/eQsVBoE7W599rYkF523/d/mlzHDi21sEXSncASpQUIibE/FD8uR8T+QSZO2Ha3rh9fdWe0
sABK5Y9Vua476EikmKc8rj3g9JHxiYRMlKLaD5Ggrww6kxf0R6xYNyQbpQ3p8R5SpHD2PXGTIRvL
Ttygl2wA2CFDmcDScwBvnsccsE/DX+eUjbiJh5gLq+Yv9KkuPF2+y+P/CO+6UKOz5MWzL/4WjHAO
QNGoXviRBXR6Sgf0ENHxBJIkCcjUwn+DQExR8XTqAj1RxlRKGhNKBI/XKTupFQwdCj85SnZTWi1Z
aapFWpFc/RJQOkp5Cq8FydYk+rUDCdqxMjtFlwY+lmLh6E9EDD62HudacNh6pScDMHxjrJdT5X6z
E3sAOCTVj5irugvrzqghlMVSRZul0+bIHka0fmCobgCG2jMlN9uIsiFIZWFu84EAo3FDAtFLN9iu
cnqEOgYnHDyibjw469Xjg9AHmS/D5trG+PQOdsnVAzS7byN9SwhHM6lcJVqRyfKzAdpp4LKlV8au
cpdzC1L4WN93dUkB7wLvSDrLlpEjkNfR/y2G6cdwTc6V2T9g400f7VyPigJZ6iUL2MQOoAUQ4fnp
O6MWLdInePKOCl6JOanfcp3xYGbGpjOrAzG7uJpVH3lTwxd7KY9ztJDwEmR0i/kWpdRSrMknw8ht
HDEhI+c8qQ0eQJ3Hj+2jmL3XZmU4nB28PfwwBGTt2RkJ+JCGpyYIeeNtMgZc/Kh6UzhBrtt60Khl
lnRbp3DYxXF33HWggfg8N4+RrGtXpZWcy4XF7QGDjYsaZKdYswWcbfaOwBtaRlsjyXgII/KYgKBW
D+XmCOtW2eCpYtwMixJVG3eJBArD2WhQnNwowFGlxq7QjILLCDjGHVht2cKFtnf3K3VWCgX6zB6F
nruIF0+Doi0F6usp2bpdEXMaJVr8wX8vYb34JpxtZeHz7DxXd/39EIBzT/Jdiuy0PMmrw0vJtFyA
UpGpJ5BtoZOVI6nzGNcpXmoXWwj0vO/reqXQGKGMBxv6/JZQv9aXNi0RmHOEK6ArukzC2Kl4cMyv
9Ccw7AX19AlryYVgK7D6illmgaW2/6RJ/ZnHV1fE+goQ5J13o+OhT3YIfSpBaIolwSRkdiNlk3X8
0NfJWTL43QmA8tazM39DdB37yZyGxO2eFWvHJU7l2UrsvIKRlhJZon4aXgG/mcfW/DVIFeaeJVOG
eAGgC5DPq6x5VXfQ2ondjea4Pft0CPmuPyaCVabT4w3SYN51sS25mI4OqGM8/6STrfgWmeh+eRQp
ncfRAIhB4cPFPek1oXBWS97ubKirDvH9b5GGky2StpqZsYuthvwQHl8f3bBce3nyL9x42vT3JD2r
MJKRohA0j6yeugaGRO1tF+QDguXTRAJM7RIqTJUluEv6ABL54iGDurnizT21O7P6/BIXBhOqpAN4
p2fEdr0wm72AcX/fusAf6XZ7761MrsJHkUoj/gJMGiqepz8oKUzW87MstB32SUv7pGyKL8zWSW9A
pZpvUPWgH4FvGbV82niDtbBaRA5ZhYf0GbjyC5ZkqBbyimGLRwlq2k1oQbZP4oPiXGwTIwTtbqZi
/Ep8wVS0XfIHj0ikh8GK1bulFUbw0hR0wkweX8A4hE1qv4q54W82q9OwiiTlP+kvml9brsv6Ja6T
GMlg0rkS0J8vEeRfHyVHn2SbP8GyjwOsW7gpay/57JpvwrWzIEsl44Akth8noS5tH13c7WEZLfaR
aleOPh68AHmr5/7ISoLyTRWmX2ksgkyKew6hs5TxcstHXH3c07uNbONdMCajZPybufgaJpJ3NYSM
nnvJSzT9kSWtdreUuV+4jnEUiyJglhC23ug3b1LeiGAkGTZrIvhmJYNQCgnf2e7Jq50GkTnvD7qh
m3DPlj3O6KCXyPp54yGD4PEOgYOGzQL6Trz3NEKD7Qp0Usv+ObR9cEtr6qoeA88ulKISLCw52DwA
DjoQWYDrhjmaubUAJDFpkFC4xHXYQopyfuxKN9+Juo/biSFE/ZdIS8oCOhfXf69CqmgT571CJS1r
K/i4dGV3azDRF7SXsFg5vVaT8u48QqR0VEa3vu2GkytbwFcN8/7qWwM/rXpP3/L1kV/EAdJr9bK8
kGOqA7l5jkyz2RSTp/PJ2sL0pbzy09qBDRZgn85iIGnUXfp1Jc+CSRwGSzZSxxF/oC8AKrBC73Jf
nLfuQE9FOl/lx6Xxi1lhwF0BNQQZudZuYBU+j+IrjvnpAaI6fbdMPddSEHxeCBIKBcWItt+3piKa
yy564D851pLiI0lfsabvAlQPi5f7goaT+1Ja0xJXMkpdsbt3pF6Tfv54GU5QHLQNTCXSctEOpMdU
VKv1AKaLlt3jwLPxmQU4qNW40WO94FHS5TJqO08QWymMcKoOUTolEVse1dOpDvqRxWIFKDxSEzuD
nEE+tFziqhbt44FkwXrNXK8C0raFPh53UO5W66Je5lOu+AhKCvz4jAVmXL+fNNmFU4j6rIMZBv+z
V6RN2IVqmFcCkXeBikX/h6GqHSDZ9U4Y+NMM+fjeGDZI94zPMcfZ2bmouc5Ti+kCNFMiMb6+w1pQ
93zjhZlPY45FrIatCk5iDfoJ1UXZ52Jz0aP3DJ4Tt9wjDYJ+5tNGPkmDcLbyKrmX1CaeYQ4zZRhF
HtffnQYobBF/Mgznxh31raLJ+hP2ozihWZpkz4vdKFHRd7RqF/VlTXhHhg+8RVaO9T+Wq/DRka58
C4+43Lty+Z4M2gWj5DyO3XVSFTrp36vh6Z66YBPvHEM7bTGoX9cU6pV/eqKV7AnGc6VZyPKGh15u
zKFYZnE1WE7Ibcl9jHOIdLlKW19/IOKuqNFrI2+Jla5Z4cXXlitKniLPjKMwEs1eXJZL0/qv6rtJ
JO1lbX9d7HPJYwoqYqgihwVdAAjwmc4Lju16UmytkHG9UDhhip8FJBTpXIY6rd8NtFf6x7uOoU1y
UTBvD+Rj3nowsWd7sea/OuJyTTzwX414PU+UPDnUQI+J28dkJE4KD5FjElhECe5I5KCpMMeVYDz0
jDBxmjj44m547XznmCZKNN1dhwM+nUF39OWikC/NOrclefKJN4pYPFQzHqX7JDQLPg5MzS/OxKfA
FGRQTwA4ARK2/lAiyXrEmj3Umbkjy5DWrzucgCOxqCjzuXEGBEpz1ruk/02dT1nREiSvbs72IeaA
wqbZDXbbZfOCF56PNhTTopCQGTwHKNP1CqSLPiPex16GHS8GV4aC3Yq44oS9xgr1f5QTnKWI5dsU
fGPR33QKFFFGx8+LM0jEfMUg/ycFGbJ/83sxzHO2723qqhDi8nmL96DtFetRWjw1cuxGi6W9HaF3
nObMTeBhQF30AwutXakr4GT/0a/nHq5dfIzgZUF+ugQj5EUoZC/WDqgRuamFR2CN8CEZg2DXyh8d
zX0JuBHI5HQfAb0FqCDQM/H/UkWWyKOrEeBWmTEY26J70a1LqDJY4+RPx3sIk1kOl0OxGlA40qbm
wBqQTEiU4MlmT4h4Gw2Uw5D/Sbl5jU5+VE2AMRVc+QXrcP9y2ofC9+joK381jXXOzDMbkpLJKTYd
2M4M5U5djNAQMrSXPlXBramAF5u+7upTY8ng8gM5mYpacuW8qLIkn+nqVWf5c4GrI+HV1EhxmswD
Gj8oMCKJkMqxVFBhu2UDgsFeOsnqROO3NxOcOlwB6c3imKO895vjuzOyIJauBP57AP0UagUpthtj
t+GCxgNK/ifFHOsFJVHlpYqu5KDHdbmpqYx1lc4POt7AI48vX4FPY1yu5UOLoVlr2haAMhK6j8U0
nZ5HH7IoPdc0aUFy4IoZzrqho4TWq5FCOin2IginsSVCDwsDW7j7TrNlvx39c3VPmmozAtinloi5
9Z9vC/Dq7BRqPbQeBfmLpJWZx8Acw1EWS8jBt2FA0LZVQmlALbn66HA//bxlG2h5mmZAOe8XdGqI
sScN1FIc9tPAD+RUdFA25n3MKmQNCNge33pncklfwce8fuAe2BUhTY4pu4uvn5fg2X0WK2at3FVc
TrjRAn9w45upnD3BrCT/BaCGxZ3cPaV69liGe8zD1PmlE5PnvMmhtsppZOEz6L50tMOg49vDlK7h
5wUXPHnbeZtxAbO1DQWpeun8in6lYt77grp4uxfA1GMssXTwdIz68wDQj34lWprBwxtpRpL3Msvw
n0Kw984OHHE/W7uGeDJHhImTruOiqSkVq3YhuFcPRB5CmlgtoRBD+i1N3iLwNSL/43t2bFzYPq2z
0IFsBL0VZ/JGPAE+GpD2FoF66L869hxetSP7m8K8epcx8lKLH5/IcOVaI53kbEMdKrjoignpQuV7
FzUG51FF+JPIqiHj7yU+qqORudsNw0/fbX7eL+edkvaodGzDWV5kPsd4POWWu4g0X9IEzC09oWlt
D7hszRnIXlVEQ/mb4pUfQPeVrE0iYsYLnLKEL/ez76vU6ZQ8xnIflpn3Furx+IjwjEGXIW+YpULO
8jQfiF448D65rmlysDGiteFvBQcuumN+1WVF+LRJx/ruzVRhVX3do4gd9FLQaefAv6PQnOMpuVT6
1+KTAWjwdtp6/COloryVS4CoTuFFkJ3V5+0CA1JWuyDNjiQzfizGQUGOJc9jTDDaQGy1iUlUUR/u
+g2IDEgMgbWA00fGkbfKfmjDWKvooeq50K4j/U6ymWNwJWKi9LusY0/Dh7CykXwTRGPLGROZHLTS
imUZRLmH4s1wgojk5AiJKO7FppLaUPp3vruT7ih1feTMrIglWZrx6Po4NjZ0EvKBt1FGs8TJW0aG
j8kQ+2/SrczD59ZzVtVMOzWtik4GoVaIk3Ep/6lP7dvQxGsZSb7mNGxpiczDJlW46FmubRz95lE/
mKE3w+T9IpFNB56SAlcm0ce1pkjKLA1d+kmnrY/0WisZzI4OTEgcaO+N/KKu276dctTRoQfEPm+m
gqssE2Xb1hNzrHNtb5lsnrunt68Nr1neYxMq0TBH9DBZz7C5TKyD5J0WYzNKOUqjDN1TgO+HCp2c
oiyrTP1iQJVpdHolW/l40/01hoavA+H/5h9DNQbufRWimtKUfd/ULCEZ9zQMx+LaDJZEb5oq19UY
xs+qDBMZyRO6/zjHHPGfbebhZeUQOyxjna75zz66NmJ5Hl7vcXdwAPKSSVbHaLUrYn3MspQJW3hV
Z7NnXZ4dX/R1XSaAoc4rd/iZQO4NtbZ6kkAxvWWH3O/OZSgN4+GzpuB8D3DvO5yYLj2j0WnSOJrl
NuL2c5YLmJed8+MZGGiOTY8mzM/8ACThNTvEh+3QhUJJNLoOovmeA9EkQxiTulWgv/viLowrauaY
mmmHmmWcoChPM1d789ncD5u99e+yvbWM1tNh20lC2qvNq8pXSwM8XRz0lutdSa/uGvVwNQ82aMfv
jA4ORVVEixMsGEJ/XMrZXLfnnqhFUfjiY9Aud078sDGgEruZD1hEpR7xkafxkYxCWqy5tgjxLk/w
/BfWtH9UA6wFuVriNpRLtQ/Pu2HPH/7Pdo9YviolEaYPwbsezE+3INVwljnsaHCqel1YJ0owqiRS
zj7DZv1hTIy+RA8+T4Dn53fDQTRQJyZy7O8YsQF7oUmeFTxI9hgafE59eTfK2HOsv+RsUnQFh767
s0scRWgUGmnuL2wjXyBrWdT2IEyvY/km+EdQjpDLKGJN9Ad6BUWJv9Er3crl2yg3Gw1mk1GBT88c
7s/oeo1ViVIZCyNNcUwyFW0XvBOhU/m5xAgDgDxwGzlMI+9MGW8spbYgAOb+bYQHY0u77x9H5RrN
+goQbp8Gl12cPnBuNHy5UNP7lXd5em55YtAlWbuzIJWZfqGfAuGSvVZDmbK1z8ZvJwFySQli2yqG
q3c62zSt7hx+u2WlGpSezC6ppFSqEU1isZM/fCJdu3JVtRyEw9rYhOZVlh3ro3zqs3PVrF5R/2CW
FI9q8bDmp1ueoUa7rMrHYLDKaZ6y0D0OQ99wLgUcfwiAiSOnUSy2ijlsHLJLMiMsgWhRr9TL4C8+
fed+PiAz+jz1yHhtae2DJr3jjqdMbHlM6/0HZk8EH0pfKnf89wGzVwVQnc9d92j5KIBTukd9SVi1
yylSKbVK772aFSiQOeJ4Qk7FyuOJAd/znYJJ9eq3aP7pIzLvPTcQ85JW415fcdkTxmo1zvxwfELf
vHaCanWGTnDWU2XWejTBlDhZ8pMNxFKvMzx2iVOXrqtoURyN9ILrg0UeCwz9Nhv82f57hcFWjW10
YonEkGi59sCnZPMp9KH6i5KqCrf1uUPNmqaP2n+MlCtwQOX2a7GG5c0hhEyu+O/JlPaOqEncMyie
+cBdtgCUBeEKf8NlakDxSxH5GNdhwLP+WIrhHo6ZHPBgoVKQTvNpy+vms8IP+KQ8oK5i/VyS17PG
001JQHkwdNHplzTjt+TvvftIx3zRoUugF2sXLdZhA/Y9JbACEiA66OZK7KRxsSDieNA8iGpKvJPt
5M32UR5QI2vkixbSQCxFFOHbFNpbZAhB+t8b3gnWoIp3u/tpitz363aQxC4GuQ0OMEHqKKuqixXm
tWeEGvy202jlcbWHaGP8D9OWFNldrvEYA9n6M86rTBNS8RUSyEbkXz4fObqvcSPcR6ET0zvmZXiS
37fo7cMJLHFRRaa8D89TchIBPyZRsRCE1JmVQCXNNcjr6lmc537bbHqT8H8spgoJtVGkQnQHZXkQ
3ct2U6lUHyDt+P3s5hy9ony7XZqyFjFrak5pgmcSwfw8xO7wzuFbIzRb10Np7ZObtig7nOqMziIu
4zCiSmdTAiZwtJ7aexHE3PypWVx6USpr372hWvk7K8eS19nlLCkRCJUjcylMuaCD75KxhOekIppU
w4ZVwjEv7tGdmJJwCtYqCrax9T2IcSyTOazhzDT97lSSvGsrWYoGO9qjgvyreKA64xRGagaZkOxE
WtzgHFz3rUOpK3YxYuwXmMne060dZnVkTDMkvcD8TDPYYAKrIsAee1WLOLCtPXm16Uo8bgcQYDcg
gqqKNXoNU4JFXPtOXQGpVN2cvLwdH1BBt4JZb58tuZagsBxGeQ+zRKVcW/8vR7N0p/DTMuUZ4jDf
D6XqaFE0cGH497NKoqcxjSYyFmcGWoFAvO24+MX26i2jPSjfhRimJku9H1fZj7ShtYrZWZin81Xw
1q1wfrNfiHsHoF+Y642H021VTccYlRtX/7GVR5N/9wK51nt+IHwi30g7qRfakACO2mA24HfKwpKa
AybiLobTxSqsWHhzpOOKH36mksYOK6YX9b8w8asZ16io97f7OBNr0RzPPTkSnlvT8wmHM1pH4mUK
4GcZx3RyhlPZ1WE74R1R+EeCAIbbNsqcgKb+KkeOl7LpEmc2ANzv/8Kfg8uFgdlWYSCqO729q6o7
2XOzpLW1uSLxQttLBIqVWINM4C8t6kzzqaeBlUwzZyf5KrJXpDLdGocM8OYfNY54/3m3k+SJ+Epn
eMITKu1xnV/J61ljwOC6kAAvtYuE+N/87EJ62ebk93jmPogPhIQhgs59tMcd9prruvR9uhdxXUBF
qslNouGqqjgFk7vdh9t9SUFA0dxss1LklDTj9HBnhLOL+imsWRpSRIWNH8EJLjJaVZmZIvxGjZn2
4OdByP4UiVHeGsHjNEMXg0vxeczIga95DG2JoaB//xYA82nUAar8fl7kVTm4aPMkNZbS8pCKAqBq
8dkQ0KrWKL+buSfu+kLn3YZ6d/D0+GWaFuxQkZ6luiOtkONE6T1lUXYxkZEQUmF5G4FmH0XQz4cL
1pKTCdxIBR3+GSW5xlYXE70LdlPrulT8HTcaw2Ju1Jk3ElMjqu4U0Afso0zYDVFyVygt1gwEsQQ0
YH7R5e92e0NROlvchFzXdRopjbuldapKlbk6IFJkKBmS+Tb4wRNppYPMDV/ZlaAS3kNlA4BU4lS9
dK1IlJV0ll1EOMp5fyyhFKNg7dlJ/Ov/2eiu9SGKD8n6B501rhzIGYS5wp24o/aXTMnj7ewnXPMf
fGcyMTQYTaH1EcFr+9bM17u+Bne65wEydNO5gyxOKOhBgGGBSgIT8OX19f5N96qOKzrEx9VgeGdh
4XI5Xf8HYru9SwZZEw50ZL2asHL0iGD+rBCgxqQERPUNTClNXSmqlUuf4q+8jDTz3RJfST3LjQcC
yaNy4QuGfpgXsAFw4AoTQIy8E6IHjUM/BkoKmFqhW5EZTJBwmKiovqxivfIbo5dckqUD0KTGAJjk
djYzRTP0bTPags/3Q8GpWlETtCGyjFpaOL08vH3+VSmZUAzeYd1LKHPhyLeut1sSqdlXW9Yn4RAu
2N18DgcbsTlwbTGkGhHpXSW2lXrX0q8DGRw0QNvY4+Is7yGjI4ThpzC42jbeHmVhYClMfhaX3MIT
ZJ5MX+KX+XOSrkiZZaAZ+Kq3j3ASqH23cuL5/iTRbKmqTlEfOiJMB4n1sSvppbjMF+bGdm1iKv1e
vOUeVa1iuPB12Q31r2+IMWwEeAVb9VGhomo4sPu+MtAQp/HGJvsUIFe11WnFY+4/SXdWwhpjx2my
SRQ6BnabmeoPXO8/T0/MM5bPtQ+4vJmYohUdXex7pgeFMwVdP9DBWu8BRTfGrzRJwsM3ftQ/1cyi
S70WX9uvzCShvjFgUZZyQwJHL7sprzwxpJE5y5lUKA2LEpagqbGS+trKRrJ7WaiP/zzWle0TAC60
qUg3TpwwSlNmK6UwPwwO8XHGbHTrncipdfv+/NAgQ/rowSWbRSVoQJWcozPD9Qffh6HZi3HzOliC
8cpV7mnmDktZlau0C47B/gN7mWLH6rLSjLWGht7uuGr/IyI1/uZoG/ViQJDZHc3uzFJE6Jm8uCDW
CpvYGkNUaU6m8KHzgjbxdvv1Vanggsmqbs2mA2cRZlGttoCZH9XzFL6t+JLpOTYrUZXzjvN5/5Br
4oGzciveUa3u8P/QOFQ/RMPRVIYTtV7OStyBi8h3OyeNbXhGLgI59ZitixPdrBVadgLY53yBre3I
qtFaO2UTDcm5+hTUo/nkRrxdGRguEFpglZoxHLFEIp2r8FOkjuPr7wZlZ9ioeEZJDuQ5zP52QEsM
6vVNeRToUgfjSOWZGhRqOG3UpZjyLDBZ6q66gwZPyddXgcYLN7u9+RkqYOGnw3vVybgG1TLGgq8Q
tS8ElsspD7qNkBpM7/7YF0X3cnxQyFKbi0o3bb+Xij1OErc5ViYhpfP80UeOUyEWEbF1IwQX70bx
bYO3t9EfgauXARqzuwxb44kNpWi47YWS2uwNkkvEuwQEofNUqCJEeLQna900ydeZB3iWxAzanjuh
A8E2oWUf+scfLy8eVg6XlyuUjCyYLzKsiT56mFlhNDfOHN5speWYlH3WHQn9oWRc7i+iGeZrKe43
HAr8h2qY9nc3IUF4NgTNjh1i+AlekS0DZzFTF341a7n2YyOWCZERzWxZ3sFiced881uH5aW9aALm
YZ8IiJYobzjcUHTE3aL4PtzJAWXmbfm5lA29Mys/mPA7MdqyGWBx3CJXLABzXzg/W8TdIL85J1nI
t38xgNDKF8D1+6Vw3wfILb8ivQytcuTZ8GXL5VjiXGAaZOligiyjC1igvqdLwYR9rPyZ90Rj9lDk
N2lmlIywNnzQxv4Xc4EWBag9U0+loP3cLdiBdwR6mLicWuInKY3Zv9n9kfrZxZv4UQLH0h/wveUR
E2o54mWBCpBrWmO7vE+q+r5h7Scq7GSRqGC673+8dQdygNPcBjvL6+lfHtDj8Nwu1TEzmrb11CXI
4SLoFYsskSHWx6doTXokVuvEkGqjyhP8KmH4ZL/8fI8AxYZvlGRawVtw8CBedO9/AvhYknUlfi8G
r/GS3a1+pT065vyo7ucb+WDdWmmnxxgaxx3PjXW7EWXmbsIZ4FoPYnboaZ/HIbiurjEyVplsNcsR
tQQFbfyAfEhF5K23XW315j1WL82LCwG9Gw/+DU5q3kuG+ONNbMsI40nnDzskZcmOWOIRBr9ChU2K
fiogJYEtNeek19FKSVY7GETYsb3Pdg86nTQeO+/9xwW2zpDnXq9nOKqUaQRyY1W2OnFLKz3iQYU2
j9fQhGv2Ux/RcFpOWEpZRk3EnyeJ+NpbOf0BuMd5zqld7JsAlSrmj2sBoxK3yVKpmuRk6XLOGJgV
IQ35udqmU0fumbOo2NDkvwqgfrRRwGrYWDKoXbvpU1Es0f0vy7pyYNlr7odVj1L7PxxVIw6aw2nw
w3ZQ6+fsWYDYGW8Qjitwdxs1hxB/mQCPQPp60U1OyYpT6XFpF55A6s+bNS4oWYA1Px44ILDYl1NU
t21yeaVuxEWSt9Wu74pa/nZhUPSIx3ao/ytHUG713Vj4C8hT8hCN4rQd9E05TzVWWtPNhvDm5W0f
mtxjHb5SFGZ34jhX5NK5GDlRl89YOI48veYmoSERKXR5/Sr4lvaywXT7ofikwY4AnMIYWMWhK+8/
czuk5v6KZHeWKaNVuiLbzCz2QwDkBBWIjmsXhWag8o6KhfM6Sf7B0pP9p0tQ+l4/oqDSL2WHVX0s
lcwkHB0Tgo5MdKaZ688mkbQnJpe84IAxRPKzCdgyt/NDF7eU5/HPS1JnMRiy20VVxhEYZjIurPQF
42C6CjnmDbOUX6TzLyyldYUojuOkoePHiteKkamARjuTDsRjgs9GnnX0L4IQIUyjIwx8z32O9Eg8
SjbOinhRllxS8WYeqizs180Mv1I3I3JT+1EfAMqYeFOEEZwA7yxUIbiKGGV6C6Fl/75rf3XxKYSB
QJtk9C6sJKGlSDPw5ztuIsnvQfgV1LMyzw6hSy7i8MAVUAgiAZSaTbwh48m82gyAnltnwWCn139n
Axn49wjusce+j9DUhnF2E5KiK9lWuRIzNxcgosnJyUgltHBguQbdKEgmopuIdHpeMxDTsdVFl5ir
xlaNKAA86Lh0lLCOqjmpHnm5lZtOABV6md9v68OkKw62LOX38BGgP21H/OPt7rvmpGKg0afVcVoK
njYla4gqYRrvsHRDX3JDywY3SgylfC0wdMbwSD8WfX8l39Ck/hkucYTGuprUHL4u/Cakgr+mwv9v
Ous/n1Momxq2oE37S3r2GwF5HNJUXx8RzAnZz9l6FU//JEiOJZNT916RpD2zi5dQLh9smD0r6qeU
BMCqN+KNe2/eHkDQu7dnUiDDCG2pjDi3q1O4lm5OgrHfrMT2IDkH7WCd2G+M4KYqRWgJc+oaymEO
/6nJMAMyraJiD4QikljzgcWkl10WLYMDRg6r+rPE96SJx1066C/cbYFO0WPJ8lXzCFUGM5o7MWyQ
LGMSxjlzyU0s312owJdhbEuCOaEqdAyu2x7clwC/uDdKNA7PPeU/o3ZV6vYkAoAutfKbZlgoL6hm
j4SdUPPW0ie9wiqMqKXb9TK+B5mcs/x42zQ3dlmexiBwIY2ArA1UqJKajtmczooUp8/E5+DtOviL
h6BiKfi/AHMcQXskBcwcH2fU2UaYRpyRSZ7j8wrKS2sjkGM7vt1vcqw+utQxn9RD/dlogkb20Eb7
FA/x6cqb7jd3J+nPKQC2eQJ6VUzPWZ8y+jldvpQe6/rHXDsRjZG8xZ+iqjmWpG4qyCIRVy1VrO9U
zOxzHMWGY+7SD1wPFPX0jVVU50WM/AmXnXa42c6YdcevLckUbqGiBoqfmOyTSVajlILkwmQxP8uC
si7BcCVxoHOOUKp8J7AbLj4hTDr8ICLuoMFKEzADEe3pXhXAu20jnxOwhZ2nPnrCX5MMzUXNntj/
Vsz3T/zieFCMfoCzgmUY7phHaHm/ieM35Xfaj7RSB0a0EwBiPzbIjqdg+b8tfQKweGGK/uQ0dNii
lrmOUG/qZaW3togvtkv03AK8LqzgM6xajZXorV3sJOYkHEbuYpzKbMqG7ZzoHBzRDsFjplgok33O
86v+6erqJvQ1PsChGtSn6L2JF18lRSgG+ee4URQtXCKGA1by/pwIgsm5lzmmQLebwScQwPcaBbYL
EHH3yZvCrbfIQsAhI2L6tIsRlqaWqTSHXZl8YHpKxpyP1FGMsc8bQCjtVLinf1D2jnECAjh71ahg
J9LoQD5P5SCmwk4fGEpMGT4DI2VNKKUjK0wvmxpoBQ3D4XOGPXIhFqFo7ukxA8tTXqYpp5PTKWwi
EI2az+csEj6peM8n8cmaX7fnlRqta9VEM53C12AGW8yaEOZX6Lttnrc7N2++6nH2H2CCWfN4d4xV
58crXIXaQ7+5KBjNY/gn57gRWJDK80UdupGu+UCV0YpTc70kBVBGSqXPLLUOnv5bUmSTIRMbwr3I
u8SnPKD7B2mTxCN0dpmEhIP6fn4fx0hpYc3ZT7v2vWV1y6Tt9gLwQTsuK5bIQCa1FWajrpSVvqXx
DjzlS6CDZfZJmMSY/DV34JM5a808ROjx8L9x0hQ3BHN36dshkyA1uiiuycq6hSBxz96IEqlghHFa
vWRz0TPZD9HUyz/W2UKUPkeooohpnRv0tb+chji9C2XQlWP5ENNoi2ri4mrV9Au/A+b+qk9Z1iGL
cKyZ0iMbMWB/WMrdAz5rNiiuTogYziL0nklPsAwFX/eLfUSWWyBrBZKKFttCbgg0Uc+BqqdwJsEF
8VuMkvd4/K5P1mbh4ksfpBZ/BohMc72p9ypNuGU4LpAsI34fOGuCIoZfwkDFbHg9P98zrNZrKmT0
VbiPFKmwQK7HYAX2nJrRHcj/3mXnSNdHJqKHy2HFmjFsR2YrtNL0ZeZIl1IVmUu9IMD0PyRAak8R
lKGlH918sUre6jECUCuqFsnb76CQG+SPhLl72WMW6XoaI/RTRhgaZg5bc5/DMFOFY+8ZaTmVIQxV
jvfLK53s1wuSVG9V1t8S1L41beyhWjKbAMuUoC8Srt6Qn+ewzesDDoKvdRMlhUyM485O8OGJUvUI
7zEknPSItkkABddam7J6ehYbEH5SGDdE95L4twbCvdWit7Ng8rtpRfcp1DGZWO6wdKNvZra0KANc
0o6cNVoPmMp+CzhrYjYJLzYZHz9a3tR1RsZR8jMCith0pmBy92mcmrJc+2hhLb3AhtDjX2wR/n6B
yknqT39h5f9VyGGUfbsG1nmddh63xaaee+Hl56z5eOSh/nQNc/ZsWMZHnuigUnXvgG1oCwsw1QRD
DI7LUaNEdUvuVvTJh5VCZNDAKHVvvrXtT2e3XdXGOuXRkX0zNOWvqSesNuhZEHFzzCndawW9IxVo
Bo9M3gFLXYIljeiFVOIMxC30O+hY1DsLc4VoBCm931+89U00pZWM86sGpXgXm0gU5+nSOqXZqblv
IHPoAtR5VSaCzlBmAhWb9rhhyEWeiZ5vBv9HWid7g9WUmQJKVz72fvGSEWt9nEZP56EzMwA/85O5
oJgqEjUESIi5z6MyisLl+VhquWjPClcnJPHlQya9igjSynC+hFJ7hVbnb6vZbcKfN6CMAEro8KJt
W3B+VMI6BF8PdOvrNP4MbL9JZPkgPAr3BnZB3ifZWmvbgqW7NYo02t6XD5A96v68KOQdVgi7b4fW
2ofrzVTrWEhp4rVuKQnBkQOzSdkOfe1JtGb/cvtnJ8AY40bjPm3t3GSlV8CoY8YsmpRbxcLiebQr
kFFVLHGq065lw09hH8N6AY6DoRrXkYg7RDoMD5I/yXmzguzb1BLCWqOJXGyUhgC9sCW0tgetUVBb
z+NGKv8JbJR75gYiTEHyds+gWnKUSGlRgJz2U0MUr0ShdMSRfuo+o3MesNZ3qVl/MWqmoWI23i+z
nMIw4hqIG7E6G9eKvF5M8bsMQjVKlsu/ld3xgOC5L/4TJwZMS+uWQNA0hRCz7PoYEIGNNH0NMhxN
9G1w0HkIYCUV0aZ9JRkusUiHvqHsy119MyrjnORmaCQBs/suwj/l9moUVWZBQ06WZmpVREz50qtl
9k2QBjn2Q9XnVf2IsabkMS5JZGnAJBbl8QXFibBJ9t8WCcVEoy7y0WJmFOjA54lWwm/ezCJvVfqG
eEwp+2McCgWLbaBc97wx23gcYKN7OMdQteW22Op2C7BYENKxh8D1GGbmyb2/9yBWETUcgKHZNG3r
1vUoAq0+cabQW/f+BxzOIrpQ9CRd7oFSliwC8r6WFOQtVGLscaO/ceR4Mh6iIhDtPLN9anppG+MD
sM1qARUChQaEFj5LW40q26I1UCYaiPYdvtumIHIe8e9xi5vcxdhDtkBX/ITY3yLo0wKo5H1IRyne
1J4yZCh2U7H4fYuraicEElgK9feAruxWrhdtBHJvhgbD+0+JD3C6s657RRxfxaSAzvL+qjb0+HZU
+iQ6BIT6QBaaKStu1tP2M8wNeW5UeVXANAksUnQaa4c07MdK+DZ8RMmAY+MD9lgrSG+ytC8vOo9U
a368Zh1YC1vaC5Zj4f0UPQNd/Ipwfi5agtwm6ZR4QrUooL9nFXEtBzylLMZJZ0IYQoMfpjx1NeIH
QwLjyjOwQh0DOv77jWo5XoaZ95QSxVdRM4Q3bNp2TDjA0nmNoGp8twwXnBU3+WByEZDMy58w6Vus
k5HwEqebUq+5ZK1Cwf0iQse8bz0ml9UdhXgAbXNUxnveoAv8pDQb9UYiAVZsrOoRsCGgauOPZWRZ
pURCq6HbO8scf2F8JzioVSGdSB8mhB2/bPh54Se8k2y6IzI8DCrv1wpGt0uDL9zV0s/iRFSMpfsT
1/0XeO73wz1zWyqSLrtH2vY8dXUvTiclHRI57ficiJFObudGJBCh/p6IDbiy4dYgSDdiN83/aZIQ
fUvnE7Qunn5BXmBYh9GoidNxmE5MW8uLg/Xsix3prln6MD37qTc0eDWr5WUB2+H9NsRt4cine8GR
QGRalXav9bW+0UM92l9wqV91zkNZgiTlcnRk+w5aySpS1Q1DEvAysBx04JFnOEDtgx6HJSgRCjTx
7w9a5FKQ4JDEEu8mCVVSLGdfQDXMnMMukYqWFnNXO30jlW4P98DWDzKnlVs/XfUeoCNdojBAK4Sh
ZdERrma/drh37Mb6JAfyJ7EPEsNVtYCztaEXpExJxeCyqyg57+R7qaPQmQmz3EdKjQLxJI+QNVEY
Ri+rnU6tmvlhwf7ej8AVjTuv6+2NIbOGp2FZ0sM1Q6S5By2HycKGxmJyUrdFPaB5tPRvS0ueBtke
W+4kV4Kkzg2+oVgz/wotsMyrj4NRjNnmD6rSsrdMz3sB24nAwFTTWzeL0SytB/GzxMgoM0xCRnQ5
shiq0flno7vAE7SkvGPf5ci5Ms+Av+8xGzh7CZN/4mk96C2NC2Jzcdz9Dw7RHkfPTh0SWnX+FhQM
/Zm7MiRUJuqOeHBXjjXYDAuoRuksz4kWxlcJdgTCZWC/GJEBH4PHFH/DNze8lQjdy02qOXXt634c
RaajEZlQ6gal9+7X/Ck4PlqoKLmDybUXNXM4kkLxTmyo42xWD8vQ4HZPLlj4mEC77qXl5OlHOyXB
3L/X+BiPZ1sxTh7EhDJmCsHPrz/M6hemCztyuZp6xzmZd1ND3gKCnvHStERuzJ4wU5yv/32pO/9+
85OoksHVcO9h5XpPLqM/ww6q2Utm449OBcpArmUXLvMYrTQ3rhdFTZbU+XXPqq6nkK5oieqB7hAJ
6smkzy5Wq4ZGKbSm/1VHfS/ckCH/XiV/a+RVwq2LoKxIGfryYn9+Jb/BsMxzUAl6SdEXGQiYQWa9
g/NjHufPNW3m5LkFcJuwKSe9d+WSJ5VYEjDu31Bq2s5Uftu8JZAsTC6idyNau4bAgJEmpxNMLLmB
HP2n0rmgQ8yiHENlRWBUPFjv/Wv6PxqLYRGsa2QPSWbopgiYg2sr0gga1xYOs7b7ptl0EBqhmVfF
Xmx9VpdfZrTXiKIEfJw8i1bJlUS6YtnoXOtjTzhqf1OdlK7qxBbcqDk8Aat8nrO1tAwgMBoejiw0
p22Vhi1FYgq4O1tRoS/CtIx0vaydcaVAkSB7yEpZQ1Mn+Zt4EnQyKbEpWfQI2cM0dQJyaKOIaQYQ
bOq+ReiQpjhy8oJg6Vm/+Qq0ihhFHjCqaKvyHwPnyTDw5BCALhVZt/+gOZUS74MpZJoXeRG90S92
iHweoqzZrkERzfdDB8KXf6Npia49kPGYHtz7uY5XLnM6NF9l28ovD/d0W2XJ6nLvnkp0golOHSZL
AqNYy9IKkrJJL5FMUv8xfvemyjCKwuBAfa+g9ri20LuxKOBIuxYGXnP8e75gk0x83n9H+/Qa3BS2
Q7XzXfz2vk9tDc6BMa30Fjv9zxYmw9RPGDoHCIK+VwnsGz7MtGApfuJFKpmHMqdD8nrADcgAJG7Q
ZUhdbAk8LRCIEbzYN/5d0fpTafCotz/FazA3JryFK9MY2cLVGgwOF30ase/ekTgNgMijskhfS5Ul
87Nq8k2PXAGWzlWLVVHnHXOrM3iP67CUOshRP+EVJ8mm/eZMLswldV4pjDBcSWutuEtirytAWEfh
PXFV1e5yl9LZjLGp5XQ9vzBjC6abO2w1z4xG1F8cGqzUouOPJMT0my7IuvJc/OZmft4fC5AaiRFM
wjxIwKlzYsVCPAPAmAz9JPWZeS2huUbbbWlePVBescu4Y0oNVdG7R381v+o8rBj/2Q4ItHUFiE0O
0rRcwRbFq8/iakO20LRyaP5GOyUNd4Y8i7WsRD44rw6eR450JoHxKPtqidNzSqKtNpeWllmG3nc0
VPf2+Kynla2E3H9MXWRYkA53tSjrsy1ZYmqZxpLdxedYieRX4/QG4g1oKUP8UxjTp4pAQ+WKYbxL
N7powwGM9SowKWKfIrv6tQpY+YgCeWUGoEfMHB41+aIk8IwcR9K9XNEPr1W3S/Nj/XMmB4uvUzQr
Qv2c+NeFraO/kLc9zJmyUNzGGnT5F21sAWI01Gy6zlaovEokFJ0VTUSwbtCn01Iw0yYjNaYeCdtp
dJfsHr2AFX4arw/uBiXV0doskk9IT7kxe8zvrYNXyC0YQXZpUYTZZi64RXF8F/L3aHyF7F+x5tAP
OygOQXCHeHyXgMm0ezaLAHXOrFCnbrovhnZMX76pfXOKYoZaDBRKBmtJ4b1eA/iKXmnPLEByQnMn
OGbvn38QyKZ2+ITXLLHxxHGKUZ1U6gWjHPpQGao+BjJcPDHiAZepF3hyqsaGWJ50Cwqrkp+ob0HO
SvtHD4vPyCiEAZm9XXbkjfUvkbfJnxIhNmZHgN33TqNo/YEPiYIaBtXQTYtHYQfXNgDJsPcrD5Gt
QYQlVhcqHLDLRx/Tb0YXdcqqbUlfQc59tVVsuuv0f+smMJ+31203P8t8tMSKw3DNq2UQrEVNgbR8
YxtiW2IVPLkvFb3h4W41Nha8RfdQDmBxMuAA5aRMRA7x+GsYkJ/mxg/DtXy5kvDuL8w5Xrd9r3XD
+RFA2W5nck4qeZ0uhbS9+iZ6Zes/C0Z5NEp8YLnv/U4OlQ06DLp4yDwv0vIsnAqS73LQSizPAhou
4VJAaff/TyhulepTcrkn9qburewAeAefIfIC90csXReQqMCEf8sBclMsiExPymleCrtwf91BOrC2
Y7m/uE3jc6BOR0X+zhc4A54wp9wla45/4GllDV7eb8FkCGUbHM2hCRjKojrRz1JyEOZ7n7JbyEZ3
NiZKEhPA1i7YJpw3QXSK5hQLH3VdFuuktVHUB6+LgLNdUBsUUxYu9T15vGuQKddwCyzVTd8xirbQ
uBcU9dypQuQ8VWw6Ou8ApFRS6a/18mbZXpXHul79nZRezlwvumgDtXzpmQU2T7aFn21HXS6f/SB+
GEBhV6SQe0owXrD/n9vDVCLWonQ+TonMA0eu/DNgAlz8MudRs0RIm9o2Uzc8WHax6yBavDyfE2Ks
waV1TlJbuqR+pBN8YbPttejG2PclFrRagvzzn9tTcEhR8DMvD1cHLel/QokWnIPwLwQTxCDFHIib
Z9AWUY9WNVZcgFrTqix884uWZmXicvxGLBUtJ9heSgze/pnTUTThY3D8OOjNjxacqdrGtsRZRxaa
qWAdtFUqnIqY/8/GkJKwZgdUmUSMjZCVqYf57SaGJoq1PQ9BVCIP1uHOZAVADft3yFcb/n+G1UEv
tIxp4rcJTV+LWKoajKuIX0de0UyqJu23mKhJ2Ij+lui4yU+jHtd+mFPNBJj/sNMIjVdITmj0fCjc
i3NI0kYzJV0D6RkX0DQ4yvPDHMqWtb979rQGNC9SPO/bQDspx+0VWPLvnjfM7EHLZ45uHTxV1iib
RpRFLefWaX4cU/Of8/3cqYD3y+I48D6N80hRtsOGkitbxCrqws0dw3LUr0kgUSMbmx8IfY++hCsp
jLguKjB6FgQhNyfnprkfkLdACkm4x7JQ4Pdpqs6+JJPX6rAEz21jtpQ7RwFuCDhMzUW/Nroc/24f
0E6zO6XW111PE4EWyP/lUMqSNUE5C3fPU4AJEMWKS/CguiaZXzq3P4FEdFHhgIjNMOPkKRf6ARNr
gZOVHkoKHQSYiwB93p36U9qeYVk+bYzajhMN8tAqi+4pDD8pWb3Sbw1aSYPAxZETg11Jac7uPSxZ
f6C15zYPn/ummWjpI0OOPE3rdamZwRHzX03kNcXUuIoURee6FS9cKF/yHwSOQgGRCXK/Oe6eGFNn
HzGfTTrrT5Ix1MgB4X09CCqZMS4I/so6uji4M2JM8o3IqhTXZW2jZU/b8Gt28cVV91ctm6WKnBpA
uR3rYiOtj532x2KILyjvdzn81a0e4u0bB02qrs4ExY6IAlHBJL3k8/HDRMYjEuZisfo6d+D9nryr
SfUoI38evmmgof4TkrKOvtpiPBxAZlAD90ySSVVwtZvHL4CcD10aYjyggdWVn8UMYSH59cASnoD3
4UN6XR8TFsxAjwlAwGOysJA3rsd2xCsMgqXB8V8ukq+snjrd83TlF4jWe9SSIT2lYiWeLJ57vSKC
KcbZ/e5X2m9A7J8QO1KbYlGCsi7QeGXQ/HtYye6Cc8QiCAebKn7WG1ptmGjcGtwYOxNlBhluLCqT
RMQphSLo+W7OIHflRar6lupoASwTB9IGby4DqYZMX/zsF0FL2B/5vm0LleySjXJR7l/oj1iBnLV7
uE966RKv/YrSpNUKjOh3c/1oM57nGFAD+aGvxmBpw1JFLfDkTozK0XxGWXv/v/RFW7yKMxCn/i99
6o7lhn1gy6MzkCsQ4yHd7GvVGmnL36eHGFStiUdKb5VTd87M1W9v3W/TlZIQGdS7CZvYkD+oZzDe
Vql5Dgd71cFBoFiOOhustaDrWO/az3O8MO63buHAcvqfxIMeVF29e/tdv4rh48t4MY/dr+MfG8RV
ZtQJHCOULelXimTDhhCq7pRHde+A9Gd1KrHlLBc0+300TqwsIKVRo+BGeNpjOndt7XPyLB2pH366
ALqQ1jt4FlHLSr4jjMauZ+8QcFM5lP0JJX+3S759wcGdKjKCbtKi29LFBmp5z/rndzMJ3THZpoxn
l/iOm/qz6EQDlfXv1QZ4/JYcazjuUl51NY6+TnNKjaqkmlTFxmUDf8ctfCQu+mcJkg/4AjdOuBa0
QzfkoYajIzlgXMLWCWqDQGJ/ya//UZtQjgbeelbc3C8rAteIdLhkDcqh/8NQSlBpjo9xVkqk0qQL
4GMwTdjzhG3EKf0GpU3rucUN1eWpfrTclEebtOp6+aia6sdrG3Baxmt+HPiS/u/4HxNwnILE0YuI
WhRS21V4DlgXrJlVHIsoNbW0o407OttJkP1xrFoJ0ff8rWxlGEfRezIoQzYt0mVzJTcbSI9w4YUw
i25dk07UHbQpGnNJpku63YfHdoHYWeCpTlVTkSdKwGfQvSPJt3FEyTe4xmNUdWA31cOJqQgf4H6F
Xf1pq+fssSaSpfqXaE2cbCF3UfI6h0GDvBeAeVrA6sBKd+eke8R95EeeZ6E/JN8GFrfOgrAjCG3N
9cPBEeALElIyN0OqMitaosYfnyMBNl+SYq8FUa06OowPJe8Ipdpko035FbaLEqK6jOQVzZYrKvR9
JfV1s558d1+iXBrEa74c9Zzv+4pEnhspiEiQ2XAAj0XPBf/xTpmTxz2bou8qndGTIZrsxbsv97Jm
itO+a26FZpJCWrg7IYeRHKfsISzZTEQrv9ZDRcb0ej/r6ilqlS0R7h7aPp0LhnceVx8JsJnzkf+y
RNR0m7i2yhR6dJLq9ePeCAd2kPTzk5C5gQTMEgpE5antpKefBOM9ccj60S57CYdCbjLRh+FGInbe
FNrIR2NA5qLsSE0AOGhGC/zGYLEqqv3C8McCLw8kg3r6L2/LCd5nFLbCr/Fwz63qs1BwcifzDuaY
/MSambgxjUKiuBRRVkl1Qm9B1mFlDIbAitA7U3hHZTLBx2Vmdm/ag8N1Kp/0wBJNXH08KwlfXSZV
u5BvErqp6tRc2ccpD9oI7fZMIyyAnoQ5y3SP6W+8D2Ahx2iA8FUIwo0UkL7Hs/Tn4GYm90m5nBp5
1Fm3gDI72N/RCeBwooS7xMSAEFka71xUCXSa9LMT7AA9A13Kwl5kLu31u93dsx3R+MAsAN1K9r3u
2Tz1gYwxuVhaB0/O+GXYYEkEDfU41PtA+pMXWpe9syRECmtnHbj/hDew3LhZpBVPF0maxg6964Vg
E7U6BYFVFGjXKl2XKU4ONFMT4Zc5gCgJuZUg6V4HZd66sNNF7ZH93FUKljTjw1W0fmtB0A8I8My6
z6twtHxK4rPEq8agWNkiZl6mLjc7QLcNK22s9Ciuz/T5kVTIGMYkjuenizxGIY1w+49dD7nv1QRO
ZYvEMYX1w3W3Rp8JXZ9Vj5U/FGWgOFcW41R8WJE8yMEAAPUwYoh5v48vra+MvenyVcg6mmlafk2j
BG/jqdX0hhkg0JlmbpViI12leijKVDL3BDDuAjCi9ZzMH2gaS5AjAFgePbTlHtrJvFtFqX3xyxfJ
EG20zl7CNzlUC+ckfv062Ft3vB2jd2vWHh6vSLDA4RU3ujyenlsPNwg9//yW2JYc4nPwvWBPn4CQ
q6nlXona9GfdeGCtLtu8kOZKVpNt+glVJ95kxGw3kfmMRM/MQoQc0Nu9B6+MzFRhiHnkDh2wpm0I
gJn80NZTAGw6KYML2nL8U0BXubl6YWhUIEPyCd1OkO66UEd06Cjdq/9pv2lYY/sFxJue8nXrx5mA
52SqDRv3pgG+aWU3TDwW8VONZTtjKLCR3KtdVS7fCic/MZC7hKIS7+u8fjPmdeqfq5VI4X0CnRQV
gHleKWnJl7DUl3+4Qr4Md+AirqBN6tLRD5xyVZvvkugpB0zet7zFRU72OB3TYMuWcxasndTWoW86
SngS8NSAInphbv/mjnP1+S8C5sgPUyqIxIY8pZJ1qYvghRFf8c82fmhUp/rq6aPLntlwCIilbW8N
yzx5dHcofuIjQsT2rj/PoLBLKsS0EnStBc4lV1p+Y0MwloXoyBvUu9MOvMIZ2GQ7p2evME7uBQKm
hfmsgLIZ6n4M2HpK//YYqBoisR9Ju9ZnY5otSH9paTrtFdJGeVIWpZoKGlYUvojCOm0QELWnwu+t
ZBH9NlWsJ9qJ/xpTo7nDBBqHghUS2ma257puIJeys+Oun1fRWmr+chGqb85Oa1l5jyx3l1zdHSVn
EpIK344k1ty59YvEgW9MHSUIjRdfwLAQuI3SEBrE3BftzSxG9GrTe0p4TzlVYbbQJsaVGFUa0OHK
+/3JlTXikBp995x+qscHfIkd/B/UfxiDI2DryjJI4XbazpO9ghDDftH8G3cw+vrIZTREoDVyUZEA
s1a3czBbDc6vSDrgQAf9N4oelpLp3GEi/+UQgGOAC5jjIoG3AmO+Qyb9OTf0X6SELpbP0dFwpG0u
UQlQuW8PF8rv06FF0++cM4quE3uCQrEyNRNSWGLnjwHxdSYy5sRvy7Lqv3QBOfmug67bxLpiBbA7
UtSDO8eN6BJPRJ00KmvBvk1NxIVAdxzig17sf/0nIRpSEQVuuZj8IWG2JR9nelBFw0BCeM8C++8V
x2J/GkCPf6fAXnXmyJv6bgLl11dLlXYIl0FeOaQbyMrMEVdTXzuaTZZrVQshDi2n9TwaSK7GmmOC
WRTXNKF3V05XiNyLGn+1y6b0xbYWbNmT4Z2qkaqPzVH5xSQBQhamYoTfZXRLlD+uhG2C9x30ZoHP
zIC0RPe+TREkZc7nPxHQ9UBcF5iLkzlPWc09cJ9li1o/Bm4G+il6lSUB9I0d/67ajDGePivKkp5L
16nRfl5fqqebszxeg6H77j9ciQgyJNDAQtwpWX3cmgbaK/vlbvDnfAoHPFTRgZWGWYFLVMELfL5I
BxX1hmW19lgFKe0pXY2noQDh/RcCh2T6p6bS9ebzM0L7ZkTWYWF7kkdfhT+nOg4z2uhpm1CuXbcc
HT54siA1VSqVHXUTdbZ1Fbr8mpZczpvcCUzUbemP3nq/r1JC5rSoOHPfTazDABYCSML6jgYcYbjm
kQsJtB/Id9PA4OJPnigaIL4adoRRyOoxDv9HYFbHSgG0j9day3SORJb2DZFBMXufuqyUGusDlT8B
7QioiJY7BHL0yBYPRfVOU919IDzw2S0wnjPi1IoE/z4aPCi26+eTRogET1RM2XftFilEQ4Mi1eO1
5j989qv3pe8R3IpsrZBpHdZIod+FeBhQWW1Ji8sYUzszGjn14YCStPjaavQ15YpjBuHBEtJiVfBB
Bz7jpJmWFVxt6JaITb12V9ydJfmqUQAmuGtX/oaOirVZCtISkTwhh03zLg8lt3MlI/hDxp6wEjwJ
lvMz8qRCQu65Es3c3sD/4i0EwpsMJAZR1hxlsxxEM0SGd+VrGa37cwgG2Sd34+biIq0CHe3ilsAf
wsxvN+qdUvF8uTJS3Wv3G3qPcGURagCAd3WEfXTZe9va09W6Ei7kXCiPtpZ1mdPsc56AyG8sWWVt
HP/nO/8eqt+Kc6/++P/SOWqR022c+KxQIITb0ANXrpEH9nW72Aj3mREXjbkbgjLf7qZq6XfKJsjB
vCMH4Ixkqj5uy3oOCcqxAGghcqY842Nb+UXYSEy6QTlVaLvsFPE9//sUX1EDgdCq2EVm8YCk8+lB
oxcN0OhvxBEB+3EWBDUAD6+ksJwaJ4jIOUxWZCH94N4HkoeVgnrDPfVyyA4vzsMvsHxXNUwDGHAs
TWRxxn+yOAHO7QVgxiayGGAuzM9egIUZZGpQy04gzS/8MJNy0wvxtGHc5nOLPVnxHAmB2DtkUyo+
K52/cg03UelxWWC51XEhhczNANQvZusth5zA3rbb9+Q2I9IqwTjdGzq/HQpW3rIvOZ7Aoe5pEIdX
S9CkOB3wRbhOctvU1lEJRXRvtovLDxBzvUPxssMe4RbxSEnEmf0QZ+BBUdp2wkaARJtO7Xcsg5Lr
SkpJN3Peb/mX9L4BAdEUGW69fAHWdqwBZNMMg4n54Dc0H7Zm2AdkZEoqDNKTGRur0KDuR522vJu+
7i9WVKDTWeIZD68s3KZFscPx2vIRK2srdSN/zIRfeYQeyHJUwwc3147L6NtSBwXBXmfFTYSossKY
yeLfr8i7Dr02TpztsAPLxaURnWJS0l7P6qqC3tEFSQiPNL8AS7dXQLHnBKBWUt6csBg0U5DVQEg6
ladH/A9JdTQeaHWuSpQnXjjJLyoRkA7BIerwZOoDlMidXdzcFdECnwvwpBZXzp8PE1BhxrmeNG4w
QE+0ZOEpRYsRajvmpWuGprQbHNps53vkimDfFndL9truMNohhgZSojAZ5Kkwr4esmL32BGemvsSm
GyqECsVz2+rqiwvy6qGwt0ZQC/FXn1I1wvIliKUiiWoLLVxooKt7AtQdVDnl04FB6etJnig6JC3j
s/ENWdiosfRvH46fXVbZJ7wZ6xrlqNRoS8OJlbpUlbkiJbce+VDR6v319Lb8K7bLUUKG8xKak5ED
y6yL4IK9r3hyyM3GgZ9Sncq+aQZs5qymvKNjzACOGF06WBLlP5ejqGccHrkyB/xCvDjO8FsjN0cA
r1KbijLs3D81BuvXIwviL9kcV7hFJv2eS09Vn/JNyKXHRBPA2sgYAa8vXQmA3BA3OmahIexQC9/d
rNN3E1CqOVMIi3IxW7n1P6UUAtpyTF37oCbBfNdbz4KzYvEQgR7nis5I2whmSX4zzMSTCK/QwugZ
P0ZLSEyhcoOI0NYvYrbonoEpmas6WZfIVe3nvnvmilpwXRD9bzTrRG/Cnu2a42sozizn6OgYHUA8
Xzd9D7Uvooe89KwUVkI+78titaJodGQgtj4YXl3NlV/KFUjDp5n20iLWWmFnYyGtmQPtRwSxHdwR
cBefXCW6HLr6ZiT5qHcsW4ExZW5dyJ8poct7qmV6tK4lEh8qXcbVq8WmwxHqJCS7RaoKCTqKloCm
GBb9ij1zDsg1X2V+V6xl2gTIv5s4bwzlp6FKK4kUDuKydhmGA4VDQXvxFkBfiR2mMwnpRn3JXLsu
4FLhkOaJcKGnF9FcXd36q346S9s7zFGyssDFbpPMBb1By7N2fefyp9SV0RzT3eRYjJkh3TYVtDDL
qWUbr87MJvpwmL9cu6dQF4IFT5FX9hh/418uJdAEXXm82zJ6SAfUbyS89ix/472ReImk+O3XK1tM
bvM8uxvjeo4FXRsVJ42a1Z1PjsATmyDMbLtAvaZPbsORNzLwHJAsmi3j9PPUe0Fq2VVfUrXPNfXO
qMA8PVTJmmjzboSEzuS72PykwXWcTASFgAcxlgAPh5zX520XAMt431EuoJ9I0E/UG/rKUu4Diuus
9rU7ZZOAA/kprSxlbKkYR9xfUmodp29IDvuleXa2Ez4llrShi2mPnuedTwYDWY7zCzI72rQvfuwH
ESgQLe9DNbgSyxG31QkKkILAHIFE7bHyVu9sfd/M4l58xt8TI4RGybfgi0/Z/QjLxxzgArpRtrjE
gP9pVHly4YELVbrnRyVbr+Rmqa2fQsvSwiusaSKIUkgPYc/RR224sNmK7d6gLlMn+kizJwE4WaFz
5igAteXVR7n9gaqjloyYoYGRG7Eygr6349EUuEvOlcv/4e4It/UW/97gfygGxGZGR0LFovHCtyxu
QNz/9VIrJno0zr8tNx6UfiQWNynClFO8po/7eQ925iaexvA27eL63GZFHu4u++htQXanhddriFMn
uYhC/qHFjWMbjJrGiJhoKep1qc6EbaDzlN8I1dMVUSO26oE5W1ZK3h50Z7yMEbKsRxm7D6qT1VWm
lcsVQhG8AJU+NF6Y+AHOYLJjWZ/BNWCxJ9+RO9UWklLS33NgMoHd0RUbECnBEIeBX+FJFsvfzwlY
uYQLikbTDwyZh+JiGYih1buY//LRJu578+mgEY98irqxXjDOKnK7ik58ghfrTOhhYmFgdDwsseY3
UY43zDc9WXIIR4F/zNAYgLEIrS1qJlDn0W6NgIj1R9gYz8akFvDx69KT0CcD90WqdH0KB9MLLCjO
OV56TpiEo1i9vz2j0BnYwLP4Gdu/rQfrHPIUahEE230qwC23biIaBYzcSIaeBAJHu+1hw4oJPJZa
AOc0D5Mzy4C+xG9zKQ4pX314QLjY56JnY7MqymSg+vutQrX/GrPEKuLkfFaYjTu3/Ue+VdkEyAIM
VPqIlegy5T4IkJzhtI1CVJCllBzYvc4spjYb88PZ1Cl5aicacNrRVxwSDZvN0ptMrYigTj/CBh09
EnHMidPZdKkAfxgQz2LWt/h56V3bOixLHxWYkKiy33EyJ8F0QOMlS2HohOSuitHewFzcoAZsYvp1
bRN2B/R0RC8jam4RG9ioEsWxGQoiGnZs3kSyTNmmT+pO51t58IRfXwa2DRUg5PaNpZAlp6dSN6as
fqyxYun/d0TFF1EDd8Du/z4ZwHeKm6PllPaq7nzmc4AbBK5kGirhq92i4130UAMBA78043ADIJBn
DRGtwieVXy2ZgWt80JYUsBIl2Sp79dVt/pkDFflJKqgm9aFPVbrLIgK7/NWDlV82sx4frd3i7kl3
ceQnIiv1uz0JIfMnwblwdvPYxt1MdemphkpNhUDVe/QhNsgeZw4vbrJafnfmnmk5ong8tzEPgAt5
HhO7xkH0idzAXu1IY47rR1EHx3kFJ56OVlBVZhAd1A9z8uw0btO20E0Ao6RET+udQnZpyTpcPpeR
t+jr419kAUJTQMXUZt8DFWAM6b/DdnZwLwIl97cLIGhYi2xZ709EYvl+NdTgQn/wFestOTkPwmkh
G0ivrEPedWeHfi1y1F+5MsZxeFKnFXj9J+wy/TT5JKoiISLcte5OKhkE+l49mCsDDGQLGHI+29RE
/h4AwbOuSl+tzFTr/0lZonOKOO+Ay4Bp0IupAhTpzjNAnOqSLR/K4FwHNhZ2KepqUR0OY3Ugn3XJ
CHU/SVCVzb4+g+Ar5zqJFEMchf1SRcHA48ibjQrQBz8S90FzvpUdLDVC3auqvJMYadJ5Rdcgd5EP
Xe5UmQRkKxZ0gEEYTJEIyqdyYywRZDsSkrcEu957d5g5sGcqt+N2g581ODC76cYkjH4MDtJ4kJGM
VDhBnq/wcY1xMEXnQ0lwE8/Ke7/kuYtgFrXCaOML/sT9+h+HC7E+3Sj9beaUsJ0ST4itTdYuAqbX
D0ba7A+Yr/RxAb7y/ArOa46FXbHm68MpSMwdfDtHHzA61Ug65S0nrNZ/lNHfuljtd8gUo3yOE0+x
LatF+/kut7K77uwuN2hBtAfRRPCorQNPXVWOEkCog5PUO0XjgT6JIM5Nndmf/l+59ANwhJhXnSl9
U0Z432Ks32it27T+vkwitR5n4LEt9P6JwAcEfBRC2YlpvB0eInLfCJ/ztNXg1Fv7hve0vKYTohUG
j0EjmE8JvbzCKWaWBcbXCliZGBwvFDoPCNkyoiICvMMZRQbmPK8pIyEFr4O4FF2t+rtPI50GwRu5
WS4xxGPUk8Kw0Ywj82+SLkenVF4Ep1RgFJ2OC465C5QJCGIYSJVxalN0Iw/iMqNToSmrHaY+n0hu
HU97oFAXbK9d0wMA4erFYyk+ZbjyCH9nod07YLiOHyBna3KHEsBdw2HRtOQecIFVmdBGmPFjOCZ4
FWynSfl/ZauWqK+oJJ6nQxWkvBucFnsAlnJ5reHewQI9eJiwfRCBTmy8eyrPxvXn49HLQ4Ixy4Ye
rI1bIsxHgyZNVh3e/9P4ZO4CERA7b+fgbJmX/enyvXPOhNMkH+Brr+yhHohTEoR2nBk74YhDeBht
e2WpBtHHSrVi2kah6qTWfj/jCs2sQ/4qbSrpjvbeWOXBHSuySfPHpCuBGj+DmttmUlUglyLZCEI0
b5HCFTER8ZeSiDbvhPt/5Yng8IlAKCCAKvK1zTwhDChbcxKBf/XmOtFjwF1++l+887cqTAvkMRNz
bVM4Xta38ifC17ZvteHhry4K/dL61rfZJwqRIrjbALVWZEBOPrUv2J19dcBIc+gt6XpmsvI3mVk2
bvzDzavz9bcb4jmZLiwIqyj1cAdUib2G9TVfrUJqCpqkG4STH0ch2nY7wlya4zceiR93ricibtZz
Z85ujqxrgV4lFLxkpGni/+l+ctH5R1S2FvlTrC9fQUDPnsETeql71M1dNo6kZ4J3pX8977LHyHgn
aplIkAdw/OZ8QUjMiPaunbK5ziWs5h24rD3Urg7+m7xJ0S+D4/JZr+wmEiG1MWIUBCXd6EwPzBa7
NIJthk6poOlGqoo/QkwaA+Mqb/7z9zCT7R6mDd2lvfJr0trhPM34n/BKw/iWOJfRn0SgNuzs5gQP
4hM5kWui8qoN8sZISqwR3UObndgb4C7hWbjU1qsetnohC8BZ4GXX/MRo9PpMyB7iP0AeDraag77g
fOe8nckS4/zn/0NkRu8PIw5zGiwHJgDV1YQjlJ3+7avMlaAYKSZcT8/Ug2pQ2XZ8ibCnzcXtIc4E
/evxPi7Cjsa6zUCEVOZRdmJlmAktU+IBeX+MWUASxSRly7KevbnE9SlbzlD1ikyFR73hnqBPx+be
iqc8Oz297UULhjtqz4Qnn2ZqmLmGpyGp2Aau1kTa9R6KybPhkWG0mcdQ9pG8Nl5V5BZyIQkYnZdy
DwZpcvsk6ugkjUYD+wulw2XIW/ocQuhDRUnPkvU9L2EC+MKGEB8+DwWf+pr2PDk53+TgTMh7kZlq
VCFxkqszSRQ4SBSChe4zmfGyy83zZHebBlZ13rTBAwpAX++xWaI6Pqcb4lNtajLPnxLbSedxFUpT
R1BmPtdtCswXJFpd4xaV5qMP5AoERrhJINa8BL22yRvVt8welz6S5YCcC0d89neMKnDOh1+6UUq2
WOnc40IiyzkE4S3hmMgnR23a8P8HFMpojMLoG/oM8hNSTOYbBI4DSlw4+LtaOKKQNoXrXfutxKnA
0O0Fa/BN+2k12srLpe51I+7GKTYXIdH/P2QNWRA3dO5SjYr9OmbBXfEy6SiQ84dG9p9OEeFLHBQ5
TpEJNZYp/HsJjVyeSFdTwmOBnB7xwtO8PElWnpzSUihq4G/O+6zBHkx3hp35hT1XzAFIepk9RRnp
sYy9FNTWJQ9s8/SMOnrU4capxiSNypUzPTaTroNXdcyD1C10m2xF/Eeq8C7+uCWZJG9kXag+QAX7
5gVP1d9RVg98iHtFKIf9+QSZBxQSaYfRA7VCKcP2PQosQzsuzmS+Xxt7vt2/QXK/JlbknTYv0/GQ
JfGf4RetRTLlNdHzoLUgu8PhvG3bKq7IrtKG0ny3TPfxmOK1X0zo28q8ybfVAmb1iY9yfXbCsA5B
JhKiHyG5/rQYa4jmEaMpAVuOtTWlN6SkFVa/8xaXwjULS94f58AjjTWFVBO/d8aO2j0M2rBZebBQ
Z999O5IZHuq2oYWU/C10yI05BXyj1VpjnUgaLzLg+aSzjLKi8cF61zBApyRz8C7bHdtITJ0X5F4E
FtLNL0+Q4ovzd0e49UgYF+v6Fkc6lmBYqsSctBoK427tZKHgFAVrHssEdsx0uDNptMJyIuwycZV8
c5sWPymc2Pymt6q9leWKd4ZLeQScre5FT3G91TPo7hdqLkBSkMVBYdhEMri99+rBZ5ECCWGghnfp
nS05qDpSyp9Oyp52Yov1FGYIW65X2ZB58wSYZcgsAFtGh6/3WIrnwOk9YkBaCt082iWvWV6egmUX
1Urdx55VnFeQ8+wiLSutOGl6lRFeHPY6ME6BBlP4j2sfaiqsD4PuAt6zTsKzHqPHEFPjSgM4RCKq
oK8nCIgXpatOWR/2ZNyADZnXoOl2EjipgfQPggZCJUNmVBuSXeWJWMk98x9dnbEDJOaqFMpeUWec
NMx8Z/8Q9llOBZYLbu+5zbKvzinf3OPgDe5MhaiL4dU/ka/3Ro+phwoY8bfGNlV5+a9ut+fgNm3I
BHyrrJK5gXD3x/58Bpn25yDYHAH0focM/SxXRNombq5AMumSrSEGbXmiOXETivYbIrn4H7+R7Dwk
qfIZi1yRA1mhTqZ/u/O60ln2noxrMPWe/AmV0PXnvFSNIJoqLhNiDWgRK5FZE2hb+UK6GtJVGbBO
yMBxOFgpE41wicHiKxJ5aHcG7P3SWKz5q4C6lokrVUKe59CMJAMlFufSi88Qddh4/up9ywknyTWx
LYYh4U/SweUjDjcHXLeVB8PrcothmAdXtorXjG9btK+joUpr+fR86khydZ0V1Xs1IL7uxMAPO5cf
V/AdYjWO7J+YCHGFydUFdQnUBY4cndIUPtAW41sbGd4sW1dLL0CrXExFRj5UinFMStCkIsotVgNf
jot1lErBjWA2iO9kPBi+z7IkPBoXC093IbwJklDAkO3Ievu6LeEMnDvhZKSTJ8Nh+AoUYoyNN6ts
CLkZohGUfJ4Z256umb76bScZmFChGOiEkArhQ2WuMK2clpXzhGwJ4rVqqCdCk/AY+l6fQ7KA96Jg
ZTbzVf1UBrx8w2R9VTDiMDN+NF4eDEMMNf36B4Rz7WTiK3bO3xe/NT5bfrQaW2sIUCLLS1Pqp5vB
fh9eAJtnYmUhkgB5oE7TZVvZUE2uJ3qDLoKLnoJX4RC1P4g26CHnsdyYEtXawluRqnKZiXC+92aY
dyzLxr1kR2HRs1vnggVc/rHpIk6rjLb9UYbHLbXYLwdrPdEq0LWW+ZLKvHk2Ko7U2zJmL+5kB2Kx
23NUbiKMSGA9IHEA3gVEfG4mo/cJfPi0eeA3KHQBQZ5ckCgMlVZXmhTPfxhd4HQkyE7Riwktxz3y
2PtWqCteHo1Kjsaxlibk9SsB+rX+0d59JirujbkM85ojnqg/EARgWR8g13gqPG25kxKUIRqy9V9C
Pke1D78JdmN+ErIV6DbVidDuv+1N/uParQswyntLGBixVEjrF2DCgfdh/TKm16XNEN3BLMR3NCYR
1l3kSYBFLK5EiuZ/gU4A3AnaHGVxHoz8k58yqlnZQ+lhrUBmCrYadjTFso1vFhQm5wEKWNIU+SAr
MXwuEWsE5RVWDU57+5azLh3au+a1+SdMY94Rxew2xGpD1IgcBJR0LPwAWjiGmMfDmBDL81HwV86+
Z7mnsRTkIIYNewq56hhX3wXoT/oYCZPDPjub4f5T7CJTqkAfauy7/588xt3AHwIaVhWJXLPUvR4f
FrzCogLAUDnJeYwpXC4jevMWGbLXgN9bHT/99ADMtax/ZoxWEzh7u9PjZDt/09K1xHuc41CqE3QP
LpO+hFsVm2mu4ygfYBaEOhfkF+nDbpO5Pyl3SadXa5DiRM1FQWvdmqJKSYL4WYj7RfcdFJ/iXaBt
aKP3m+Z5q6Dj+HNpQHxxpN3yLeKLDavvl/c0Ri1EaF5Y9A9SYYkCLLhytj519z2hfmeVaz5NLPOG
hkuN1DbQHL+GHkJX8/JiV7VQvy/iTtly9yu0rwSDqG3WC8uOB5eCsj5s7cfN5RwkeocuWzLRpEu8
RmpXTsHdJCXJ6lgAqwVhmFBpwY2pSDINCfDOEoia2v8aGbgYVGmOSNtass8nnf1Tld7o1N9sJnzN
+yPU61cc8kdHgWDgBacB+IyGzJz6PCiRNXfP/YxmEiQoCLRY/Kywn6hSpuGp9P/PbUoBOsnEfECH
JTY3ChQpJk5wZDGunHXVx7JLk97/XQsExo5XSySRtWra7mpwZbHa+lBtBz8jhwkCq825KAFKFOWs
XY/ox1ZPlH4v152UESUVeGflzOacS/7nSE9+JArrUJIFvsrNbIrRiA33E4E37dEbwfqdmAFdgsnU
CcSUPvPrV6sC1HtGy5nulzqYrMtkbCUvYxP6ZayEstg2/AONdcbFblNb7uUezhXBJg1t51bG0DrJ
R+LT+uI8fqxuK7pDW0Tl70e5HOhj2XPpxV8Wm7mYdkmbt5RfRmTc3qJ+W8d48b/UZiv1DTi3VySJ
ZtRj9TcSzvltF2Uck1Ku7X0gzVwPdjJCGKKOkJNOXgrgzShXwa9AKKiQs4lFWXtpnNjR6L0xB7DU
GEg572NrmOdQFn0GeYgz4WxQVa8oirDE38VrG+IC5RI1AHwsdzN1qNj7ctZtnbQ56em2xP5xGEqt
Y//CGo2lx1OndguCsacDXwcX2+ssjK6LY+TFSWcd2uYhpQXk9YNi7gzBXwqf8HFzDLTABI0TvMtx
MXB6Ndbw2Yg2kraF2zFVM91c9wgTbCt1bST8RiD74z6BrCXojyTADprAFv+Qi6g006EXLWzqxLwo
mdMkAB7sqDS8ExCD4ql8/QJSDZqJ6XCFazWfdGn7zZx8WOyc2aHwfuUXkotXeB0evvzYnWAfMWYC
qXocWNoE0gg/nmGtrSILIHwS+bnIV+JX3Patdq00xtGnPfxuDU6Kb1aDZz8CEEDiqb3uT0DJSwEK
WLoeq6CU6T/s6v138iLJC9nNY4ajp3ny2IuFIVcP3IVkwQhPfkdSi2ldiZfoZOuC9mSquNxCf2/8
1mfXyBlEUHY8gSh11RiROgTWz8TOJBOHtXWxTrPm4jx9rbo2ACOSvujlDhBnJ5x0Evf2NAV6vA1z
3QaBF0rcuxl+VY5D6tjfGnFhmYbtyfUVGNUxehezbXjkRBElwfKeT2K7ImtGeZNZepF08mvZjxSh
BKzJvqEBQ1L9/DuZ1FuAo3mfF7FZoL8hlQ7gkpgaaONhfJCTruOY3AL/DtuXSinrYq/aZqwX5Zdf
lkq0bbArSLWObe3V7Z/AYp0a793Nb4DFGVyzgDYmsB18VU76Qa8G0JBiZz9BcdIir+klxMu/rUYw
YwMiG3ajsl/HF5ZWcAuB+1FUXGYhnjRrmSjMCnJH6ePfncLNphKHzBS52OBEqvvtfR6SlOq4aa5s
4WPLPqL3FJHmIlhxtsmFKGgfnPHwQY6ePcBb9/H8pr84Ts8tIoLwj9OvdFr4IsUHJq2kqA+YhKMo
+7zFqDsCnnpI/X6424LHpKCi8dD4MVqENF63e7fous+iQbzTB3+wazTETviFcj4JJ6EzfGQ4k7UE
mQ+WKMRpM2eMY5/IYcyNDTlZeJT4Etqy3KVFN68rhv/6uxcKoYhfetCEnXD+GaNKiBvecEJ2LeYH
OeBf9tXi/zH4sGUomPbjIkQHFwmN+1ennIcZfEUwBY1WTgacWr/Y1HPQZ2DEHEsBGe3Db6AOq6wM
zyED1p4inhgVykpHzFmQAzF28kwBQUdjDxDysUB4ERI5iBHEKnZBtxmhu9RNh/643EcimI/7qKpv
awrC2rXZxYOlJ4KvaUWD26Y4Hz9kiIQ5kEBZRkTrk+Z5xDI9xpaH+EltOIXntdEIK0sC8kMVmjeM
+LCqGX0LMacQ7CwUSyEZWx1VHNV7dKFOqTrBTKnH5pEudBEbsNp/20lTZj86eEzdlX6CB3CqP4QG
MyqbboXwZIVGykEYyEICyPGkskcs/M/CwPtUYwQGtOT8liG1JUMi4usY6HiBN+H3TxVFFbHNIrYt
jwvpze7/VdrOJ1g27iWiiYJ0ea7ZLL6UHaTAtwjYE6d6eZGMJfD+e2tMo90OQAFL22OOszKrwIdi
PN1Io75wkRe/xZSXqAmtCXHKyaYoWnYK32TCMBkA6ghwo1VTgZMVz+g/vvPHEwbeRyiwqkElnBjc
4uuogNW2N+hrPl69P4O+6iVJXANr4URBIffS7dnQxV+GZiR6MiCSoUbAaXuv8gru3ZQQpKLpcXW/
IZq6z7HE6rN4FP481J+HKjT6SKMJMFe9SJVaEn8nG8GJzPKnQ0ItNIh7iCIJAXmeETecT7jvPz0i
ngdCaoOlZv1bFHqWmFhsdFlFXmuy7vB6ScoL33P7fKM+YOGnLUYttgTCqe+0dzB5FOS6iNPeuwn3
PuVerOj/0/go8zZN76dtWzngvJ+tfO2zAhVzn90sL7sPp9n5IeNlUdRFPlCPGECyIIn1XlaPEiTp
3YempicrGNAmbylM54Lgd49GoaMz6heLG2jS/4m1sznfr/YkJ2ydVkyXlBIlBb+YA8Nvfd/68pg6
B4v84i8RShOKAVi003BW9k5cEsx+07BeNqzZS3yiQRZH2EU/1pn27AbjEuh8Y8/oLCy7xAjKCslP
7PKHD1wQrlZJU/MlVsfkeuLULOF0FMZDecqNmb/gj9sUzxyPBxE+/hQ6/k2Y50gSFs7CES35ociG
70BKHe/qvTZWszFTW167BywzhwSOlj02ACLYwE3wZKX22qXGVpH5K0Rvo/X4drLHvVySnjlxL0dF
zlPshmifQ6Z/8GCseNoV5eq5vRZHi4FqW67Ax211hiVRmq1hG5um7S3We71HoGfs9KqSk6ed7B8F
Wm3awc5xSFTgpqu0jXtG/ns8cQWcGZoGlrOxzH74TG0P8FjxUOKPtES4E+cIltjS5iiPXhonaC/V
Zlcbkrm6zMYtyIIZray1PnytzS5uhS9A+dF7WZZ06OmD9/ErC2ec+bGc3nc2cRUbbBGmN/ZyGiY9
cf7tq6rMNDvOFrRmBMjkwG9kVzHHF5YBxETNHML4K8cfL+KdT/rV8fci4LRrSdra93PAhW4Lr+sD
ZRbH7v1mPtvq075/OalrsX7019x8/vQlQYBGpzBef2+3cc6DGceLHM+Xe58Yh31S2SsXPXOl/wVK
t+bnoJ8LolFo9BsvRcNxd/4dELIAiWGVkNMpCZMs/MsVch+e3uf1U4f281n9qg8S31EEzSEVSM53
oNaFFhX+iD9LAWIEFz6Sl5pkpTs3njFUHJykqcmflS73pQq/zM3Y9cwLwpYyQvlf1BG7VML9/zMK
O6uBeMySBZT8FeHU9M6tB14fRFBkNuCAUm7tbovTBqrmQlOXYhYFfHG8Q1BxdwydQU5hsl0ZVwnR
ZmtWls02YatMaFSh7ICNJKaUA30yBACzPOkAGGId8+zrOz3DUzjZRLTtoaOqyaJKqlzM7fXwTaXP
kPG2DklEQ0drccumo/Kob/zLbaG6mSZ8Vhe9sLA4p42ybw76EurP7yhqxhIR24wMlAYF9RWuCOV9
MKcY73aa6yGuuDUx9KkoGaq9ehaaSeGwhqWWUX4nOSFAD+mtKjW/Qy2GzbkUDUJVYP3pB/FOxKN0
LeRTyN6JgaE+fJkWznOQORwqEPUbJZk1Iv0rGSpZj82CMPS8+MpI9/JzUimeg7tPk4HxMYWUFGag
rI0o1fdT/6jH+qMdBK5udWCCYuszwfHSqSYaq1liuKEogwE/zOBi9grKPSOcoO2CC5yCJ455bRxf
Rl5oJ4rdwscMKZu58ndoW1Ox7aXyrpx4BBfPRfYM/i/X3nQUXp/nUSH8N4DFsSLSq5qnXxztF6wj
t0SH34v7ZJZFec2V6BB+oiZMakNQ7pF5qsarlpcUzuZZHNeJnTXgHNBp/pKUBht5j6KHYWXz+l4q
pBY2VxA9OVQ5eIAPfs0w4Sla3uABUUAb3bytP9m+Uz5FpB3TLAWIzXZK+q5b9TdLvnm9XyY7PH41
6WUylSNQTKu5OTDvYn/1tSwBH8LM7nA1rkMisPFXOzta+4PiEl8sPqzeM4Ys/lmopKrJhgKjwiPf
y5lhwgqJq5xCYC8mGwkogbv1bzgfnWkXQiMO8QSvx9R0lvvMOoL8K2wezgDiZUy2738uRj70iE6o
c4GThG6wKdFf+OoFblZtU+klo9rzikdNyMqyIFNMq9+7uR7a5Cxs98olBcxyr3qLhvQUkcKb4j4w
8QqJdoOl2shWei30NIQ8D1CIJrGRwTMF89bDvHlYgOLhStP/eIjuUdpb6S/zg23k77uqXhK4c6SV
/bFdVflGFKd9yK8OaxY/PHQ2IN2eLcByIRhdrJSOz8iINRPVpDOZ5WN+Gl/7gt89L3fKS0wujt9E
bnuCjzwc5qGybhdW6yqrT41YPxq2gWqB09YLJSJYWAiUlixdkoS2dBsW4ouACRYxX36TovYvvM0r
wGe3wEEgEsN56Us9LE6WFcUEE4x1LUg3VDyxnwaSWh4RCEN0+ggOweIVXtviKV4jOGJ9KNrZBYUp
yy9GRuSu48SljHkb4KJQSXzerFhgNcbJOfhqYYxTKCdZD/F2U+0+nIX8HOTUXBx3XCpCS/zcNWQw
ATPwsvk8r47Bi/kkRVgWx7UqELFLkdXsF2JPh5qH77r1XPv8w2BE1gT4VoYZYo7iexKaH8FmVbQ8
e2AaHSBwBtLIbFjTTjsAgj2GcVGl2jDS0oqFQcrC1QVD5OD8yburp+hrc6tUtbXN6pn+YUpqdLXC
osYNu3wL8j63x/5e520YCl/0A5+Dw3hg96bs8mI5YGcbSBl3NoJAlbNGB7CbCABMclXuG8rsZjSp
/et4TBBEsIMs9/wyX0dRDBLY09SgRTtcG1mUKpJ40CEBBTFRbgR+CQKXvMfapv/T9duZT6X+RVnD
zae8x7JwF3TWMEaTwhhw0fTHm7wQP03KPjrnmBKY2ZK9AyP2SyBs3S48P4bGhlXvRSOcACV1Doat
WljMX0JGBNbWZlnWxlpI/y31XbJReRmiJ83/GoGhrp0Z9DWg4+QGP1O4G2Ef8LrXao9i4chIEIpu
f/RXDybth13V2Eo2i2pE/ZHexxxMf440AA8gNYDSQwEV+in3Uj1LkMSQU565iRT6KXeIc3eqGNMU
OGBymaxammHqVQu4qAdt9PP6eQB1sHgdVL4Pt/PwMflq7jyuclg+QJ+SPoRmR7O5ytw7s9PZ3xub
7VcFtny63YK2mIYsDwjFDifVzGLZF9js7paTHMkRLNu4/6zr4zyMV3lVETl1sue2OYvEfULG5sCJ
tFjkNF0z5U+3RCohSSAJ2TN3aaFX1BHmVjo6ax5+RDDwRkTAb8BQlQObw4G0ByK1FEmMErY5O96e
pgOtVseipvpSgMq1/K83a8ZKv/iXEzEIQ6l4lczNTbqggD4fi7rbW7+xDMrXUcOplb4sJPE7GxHO
+MbVhG4VS/L0OlnXKL31TNi5I8hNrJyqD9ekszFkk28u64R/bX22ol2qdh1MIQGyqX3vdwXVorOa
UVORVpMsUxyeVEvkPvGw3stb0/wrpHpPXU641Iom6tFu+6YgNVOnEslHJ8OASrGk3aaqaBzSVBWU
+BjbI4a9K/L8D9EhZVgXpxC+wiqj+GDhHnD2md/HrAqi6KTRF8QfHcHb/Y/0tYIzWe40IycMN6Ov
laG2prn8cT+0yZEmDtAzdR0aVNMa1YJ+ChoXqxIhFraxQ3qWSQ6CawKITyg+IqWsglPpjUAt+dFz
+XqNMpeneMkZKTAFlkN4IU/HMLRY96IgzOHCf0ADOGku1Rl1dAaH9U017MD1NxGw3UsOyb+gZytt
kOyJdkNi4V03uYHOC2t8ZWXeRL/NA3dbVzRb7K8bj6srMPwreMCRUC2JlGCvZJd1p2yBFLjK5Nm8
XZT4DqSN7bdmw5PqE7zttjuYiv/zQHr3SQ1ht3nt521mg+U0Fh8PPztJX2GIvRwmoaEt5QRrHC/Q
TQMTqU40FTxbCE+Dbsj3ZrYQm4rFFQsPwRqZaT5eVFmCcCkh91O1JqurhcSo+6CT5fYyyzFRBqKw
PwYY6khxkeCy+rJWLtceAfgTP01WriBLoOpmTjpfLHi29ex6+WzFxgdMv3S6HF8SvukUOogaMsXt
Ntk/V3fAKkMFF34XOTiaNNg8mtTm0ZoM3eBAsCgTD8UKQ9OkO2TgpOVWp3/3lucXLGW4Pyqk38SY
NTjMhY139cCA1/J9LelXtUFDc7i5cX+QeE6QRKGmiSTVM0amA0TxpsbLkaSDrhy7LT1Jx/gdvwtM
nCQThvzOYJxmgnOLxspXwK5FiP731apOJddSYv05uOf2JxVyfsNFi21F7UtQPcMLxo7pNXU/aXfy
H689Ha2f7npmecAmMl0wG3sldtYADqTJyxcdfu0iEte+iiS9oh7IgIjLItPBohn5gZ3/IRuDDOa1
yudAL2TGxMmuQ58xcaXwiZX9AOnDKV3fdUt9XGFVfpzUglBouJSBI53G/T09qwCzIyZdYm1PgKIy
xwdPRR3F3GVXzQ3fzy2xmwILJXA7TM+D5xIMaIzlZ+ZUH3AVo1UbwQ5pASNGWyDmFYonNR5fJCiu
CDZa9gMVamnSRbSMqDQE6BFE4qUVxFyKjNej3agPidj9hd8XVNkkSAScaWvB8YHBOEsoDkYr32PG
4ALwOEUJ2SpgE0vv7YVj5IGH8j2zYNJcoQTjfblmupQJz3Ila9+h4ny8TQTcWcafCTpIj51DwR96
pBDOjAjaBZIo9WsCqFDhMPIwGpaV1t3dh+ebflFocOIijVV+E6QhCBh3Rng8dgy9suWaGo3jDbBd
KPUkybnpR67ZsiAFsGpvFJQ4t1hdtwOpVMf/4qeP5H73cTMZPVIYSWx3MEnzua54BKS3O9VNVHTy
4Wp5U5aXVlPWl33ePzvD0SesBXEvqnKbqOey4xVC99HczOV76kHIBZXo5RywBLcEMvSSt5UJvx08
FxCcPwAJgQ3mxcE2pMVTJIfOS35yXEZEKRbeHKPy2rv8Kohhb6p/ZDXoSVXJDhstmeXJOzJbv/mw
F/ZVl7i7ez5/lxTWol1Ejo2ThUCt+IH/zRs00I0nJ6ZWvA7KGpOteLHPuIjWaoZzssQdq/ifBQUh
mRKgsQKxH2eL8mMud5Cf39W5PMyKH72Cg/1ebBcmG0GMlHVxqQ0oqGIcddtQOExeMkengC73YOnn
Rxp4uYpDDfIMoG9zs+oIZI5wV7cgnK8cRQUvZNj5ByIuMVcF7QdKo0XKqkGmP2VaTBvaR+38npix
BshtuffWHI7AJxKf5XoMHfAMOAIOgvcAUeui+oPr4USs5KBm5bRBtwW4jxxm+oKXWH7PsdVi4Q4n
hHzDPkPwoL0nBx0h/b+2Wno+3OnYjIW9tTrktZMoPfBUfusd2c/3v++51M1JtFaQTdzGc+4f+cAu
AP3FU/Ty+IhDqYcnR/MloYQ2BYDirLb2cWGiDr7fW+zoCmn4+DzcTTlmRKn5NynDbgILXkvPl9ir
5P52YsVfRGz7E1So+OBppi3wmgZKC3iJxatjlsWt61u9MJz3yUWBPSpg3l9pj09bkO4iozaT+tHS
/luSHNTU9befLk5zf3hBUlGwgN8y4Wqw6nfYCaa2Fj3Vfe6vdfg4WlFaDrpctfIP7VXu095d8CBA
Y3EW4FnDFvdOAPIRz8OR/pKK9IyCpAnFEhBNQqM26YJDv94BGGK3HCqWr/UQGWtv1HMze5dOqORN
usE/jMpqPhV3M2Ir78sdb8OZkTfxFCUDa1I5MKL2T9PVaU9l7MTXg0qFGFykE+m/HuTCCxOj088G
xGJMoVaQ0/JXuwxrEuxhpqUiV8QzyvjD8kOsGaquHioJLWWxwqKNO0Xb9NN6Ravgn7GDdsDjVrOt
ezIgk8HCKZyl1drT124LfftFHwxjp0NBqOe8pwFARoT84AJH6fd4Iddsp2AkIgEufCh16kSH4FTh
Q5SS3pYtOuBqTqDnPRP5Cs0gwpxsBu7Xz4K3lzpSsviB8v9iqQUH7XZMx49XEeX3NwKWAH+nhYjb
wDjxG/+J84J97nESj7WQs6CZE0/SJXtDENiErCkycAbPplxuC5f4t6DfdAklC6QobUbuJhkbfJRC
ggREJ2ysQOjQIyqL1u3eopfK0o6OJE6zrRHuIYrMrebjcg49Fh4WhxPfYqiFPV4pnjxz7X7+jv5E
6ldsDYEIVvvCu+EhnPLM6idko+pW3n+bL1KEmwI3kEzG/TqWLzEgfMycTyzHkmCfNP1/FRA5LplG
RCzGw6tA9ppSs7J0e92o8a/dYVNLSrACYDl4uSYb9IwZ7ZFdfWUGYCaVed2O89ky0ggSOaL5NK54
uxOmHZ38VJdweZLwxRFaAYg90UwRswaLymR/u7VQF7IPgCp+X79UcSn2W0fmDAdre/SnEsOu99JI
yHI5OxmkKmhzXh0oG0B5PBcSlcPaZRKbNV3/r8ZZ9CKlPTvi8t3HpLCdJShM8ckD70152hgtvojb
zdamZEHKr6eLk5J2Mu9kBgAGkfY4n3nh6MOXjS6d4fhVi7MwYca9dFttkcaUjMUwvhZomLOYnAin
j9ZUZSHJmkW3MWEDflYneregoK37LaZoz4H1hFBQUcVMFvysy6oGnbi4rnw5BfGm1E2F3keuBFHB
37ttYcZ4qK2kZRw7geyRNt7PmbcaRsyLRnRJiPI/HoZqxAAJDuIBsDByV9IBUrY3pOiManGChWOZ
ACoIrjF7MoSxE2AVtVVOuJroaGnF+WGOSAr5T1qmJXMQiFIo1QlJcvPGTuHdmVmYtwiXyWbALZ5N
g/fleArQtggKIvth7Utmh8bHLV3e3vkL6JF0by3q+pnZ0/i54K7hkWrc9ztXir9x1wNjJJNNRU9v
YBB5SfU3N1tJPySoJf1bK11Ih1CNistxw4lkpw81NBLAbiufwhGXB2hdZOTQuowaqQapBWJBQwAh
8C10wlZEL+AUaSNw4EBwNXxwurm59S/XnQJgU4r2hif8TPpx58BU8WaES7e+Ltz+uDhlMh3xl4Pe
6Sae9Psj9OOsCq87UUkUNikFgYJt9l2r/D+He36pqPYuDbLGZKghiTCFPR6MoKzddNwgomG9D5y2
PX1uRwvJlOp24oot7+PvJ+7u1CtzSfvh/UTI0IQnIZqi5vtOfegKli/oBCYdRYY6cePLOomTOLzN
VF/DCAEQ210aMuWj86R/l7CT1SgMjD+F7l3pENY2uyoY4V8aZC9WaCSBKZfk12zspPdU5tER7Cxe
7NkCYWlg1JRM8gmtaJNajZU4+a2Fz2oZT2182Np9PriOltLSMSG+umnoSoJ7mTiDXStpdOiQrykD
aRGKxOG3jTU7wg25qer05Br7NGTA/vNnguAFpvk2e/B0csAkD5B65Pm9yViw4W60tONZXEUF+3ME
epslKGj+6iOPHHNzH1DJQQQ1o4qQi4BTmEiAGs0a9RdOw3G+kVgfMpWXMe1Bj73i3W0qjET82N+c
A0gOQfDaldx+vGaF0KOKLM+lUFdGiYJTaUikUV5tviei74O6oRAGSQUPSDCBy30ulKHE30gLninH
JetTb+OintvndBCZb8U6W3yfDYynSK/nFRUmHfnL4AvEd7BLEYb0cj8lFkDL2Z5hsNKbngIvUKTq
eArpr28xQzA6DxTZA66EJ/N9HNwR6JZkwJPYswuQCLDQ/KipogAVQsXz13ofi6AoBwgtl3h4YkmS
HXOfZ1s9hxWRczDRpDCY8YpX2SJtI46Dqk2hxgo26vvAXMJ1lvSwosk8CFMMtxHdNNf28tr8b2pD
EAyFDtm4NzzostxOtMDBI/4mG7ycIi5cwlIUhJY2+Ho1bwZqZBtAkA0m9jN54gaTFt1PlRd2D5a8
yt1VFPtVV473ByhcP73qv+utW+qynKoHrhCNm0uaYRADdlXSZd6t227NtyyuKqdhAY7PVart54b2
MZJ91KHpq7YI3yKletVl2w/AG8UMbJkDzGJK72eSKh8cJNVA7hLwDzqrjT50oCMgKHoAXUQUezLx
i58ijfGgM6duKDiu+di80tR/c1zrbWzbyTMi7e2wYfuk3kvlW4F9ttyr7XoGrHXLwqbaSrqMfeO1
gtRAgNHXlEyfCsfuN9u7Jxh3pM2RQGhvPRSaEldrmXd172eJOSXk00MVdjnWtsHphp2vG3kdlfLy
hwNqHO7CBKZ6y7ey87ajrQe/5Nqq6iOeV1wqQlcaCEbEiZMiJCg929GOvYDPrP9EpuItpZk9/ED+
s6Xw0Ht4Nl9YkWeDfYQTBGmwqrjiuCP3kZ4SDZfUkIftbSfLHL1B5qpHUgptaITo7UqXTHb6Avgp
dpDLx6N92LZLlV2tEUdQ2jDKP7JoaFwu6+FBGHu422iyJVXQpsyptIH4FgQilywLpm7drBlnD+Lh
GNgFc85RZ54W6uDzNXqSStb1NvN0GQQSp9SbCMQ+6Wx/abaHK33zi3XH7X6/8ZWln+NHM1tS1Y4u
kPoBW9p+PDLddQzeekvh0BwEwf5WZD0xL7p89urkTD567ejvgqsPG4ShbAf+zI9uwO+y8kiRSx2c
kqMy/QFIMWyNcIEug/G+Kf+sA10o+RttQJ5EG+dv0TyG2TnDKrqQLZ7uSKEUsbPB8ffje4vOKzD3
wUXUy3KEtcYdSXXGw2/Vji4zjkXyjF1xeKYgYimiyUM9fq/WtE2e/BmRM0IjbNjt20CAoc77frla
SgsTqryTOg1vHbUjezjjcI6chvj5Q1nis7Yruw8d+7e2SeYYBP2QFX2V6Y3LnSMv7B7dUg08ZsFu
cZYt91UUGo2i70CphMoOX8hvWEBqi79EsC8Z5YRwXfm0qQifszsBtLX+zIBI6OdMNoR5B0op23Zj
8oz3ygWnP8xRL4mMtBJVc4L9sRaFCXAfKWQ6SCWmeOdQ+n+ou8i80Czeb4Si+MlpaN3phbEodYgn
mTVZq2qA1DcfhC4lN+889cjRWKn5ZvK4olMfIY1TaNMeP8xqbrtlJ44N7ble3m7QnevAVvkMQH57
VDn+VWRf/MJztui/JkDeYGKTp43cJgqqALVwJ+Flil8hjVT4/P9Pkmtl58KzXea678SaDlgCjnyh
6MSBRooJbyCCpodCkUoifOVikOXVQz9PsAd3fLooXdkg4161q+AKNNA7WAfwE7TCJiG+AmKfGw66
Yq8XMUoX+NhHDN/wMmI+PSZ09vZCSsibTTbDESPXb+ymSQ1bfm/d9hy1d2GaMkDSAAOegLWXjS91
p52qZkwm1UuJoueRSi+2z6tp/V8xgprSD+dWHEyTqDC+2WubusnQZLSv05yb2ixL5xJfcUgATKTX
1xcq9eOksY440kZyqIEDJYtqnyBEXTepzJ9on9AwsUIHww5VDP92Upd/3xLsYDz+ig6xuJvsnP9o
vEQpxUJ0SKJD3Uh/tNBxXZgXb+PrM/S8F7+4F1Q9UDdAP4eWls9ud4+/7aaTWiwmpiIKazPlw1+j
Qc3rWOkVhA5i2aUB4ENxdT0NvOLYsL4E9yNI04KaWZkjd6QVRBrpwz9G1fMl2gI0voYKBue8rCRY
GPguVw6LV8xYYkyWPkZomaTCiiJkSxgHj33AgyZzTSRZm5oB9QhHzVnM6OdaHpw2fu+Q791VgPCw
JCEscN8RQGki2RAV91FZTlGfMo8EbipX/dnibWjxuabTsivpfA4fBGa5xXczv8gr+TcLZMKe/5L4
WSEMfZPd7GSuNhTYXY01PY17pqB+OaNqChTCct4aTT6dA4r9LPZLucyNx20KuoHEA3Acpi/s5jFs
AJLsC06NOLWab17Vh/Aa4nhf5U7K2P07jBIocrYcPg4E0+K+mpwFrAhvyQpTaG1fDMUxuSNZkAuV
J74/ArMPyUpA5sAFwidQgty4a1tmufqpok/pJiCjOYUq7Ll4DpbmKMSgJMQvCYEHtwbHr+zv6Ttk
wYi0yRYpx/PVkx6qsW8CfylAbIl+8itL49yZ+HL0qmwK/l9D9111MLfKTmwJaXSoxu/VRkbwWOoX
CgbBq7UlKdKW3yYuWxTRBzWbEiNyzrMD7DDg6wCH+ZFfRoueRzkjxNuBKw2WBtPN4xMUNGY2UtEN
Y2e5ezc4MLy+c+QZTiSvxNNvJKIFFE3uh8xjXQhs2Po4p5QT7+FtXZ+3nTERJOl4C7np3BDY69Rq
5uo7JjdfboLiF1BJ+HWmFyWEolpcrr2CK/0ZeEt3hpcnKXombnzOYDbcwQoAYZK/P87gRic7CWN3
hPX5xUhC/6a6nVzcJIzqKuYkGTstt/IL51G9Ygfcg+/7gdyHTrsnot0dcY5umdphY4skX1RwdYpJ
tGV4sj63wzfcWuFUsSSKJe6o74oWkfPR9GkRHClQVyBCiRICWzQeOscXQnoIyPtWfmrujgiXqglb
4cEnaB9ePD/j4BPZgpfEtgyTJNMgbeuRLXbsIWjzNHsNqPPz1kIIMxqAHjSSCgjgwvt/hvnJQTZs
yLxPwyur/X+DXKQeOYzUxCLXSCcrQYdCnaNXVV2WNJwcOLkrks+piR1EEtPRVWXiTfAaXS7zoEdc
Mj4OOvhPsRVFjdCQwl/QAxysa+KdL2VfIgvj48Mi7EQFYmBigx6Xg8TE56nRl6vEtpL/nveQqxeC
ZYx1m3jAiG4XBQhWUmJwrb9cu/zu/dgBLpgl8uY7ke+D11K8XyzQopD8A44Q45ZEOK7On5bWmO1u
ETvmNMypf+V936voSsBC3d49la5yDRU1liM5t2/Q6fDaISFo1r/9o2JWG3aciZWrK8Us9pjL5fLf
A3EdMr5Z5/cnU3SbZg0cTJaf7vCiigtPNLGEyu6Zv+JuaZn6i7qzi6Zu+LyDsMktef5si+AZ60MZ
6YyBfneCGMb2givGHtdvi/3oD4OgNaFV+a4f0DDYqrG7GCP+ZeHGeg4GfVSFollikVRBjabvwwy9
z0CoyUcYa2GXtBj52/Rkg4NZhX46Py8jI3RtQpYpjUQVTB2De1wUhXuMBUmtl2ju6RwnE2VdAxHg
IZIIpOfR4rZ9Gnc1dmii51Zg57NOlpQVUbsgzlOZ7/7qUu2fGPB966WZURxVFtmVCFEY1e/hfEIw
maeCyr+FnV95HPmvFBkb88G5tjaitEPc2p6qGx8C4J8wSL8ZeguQFVGuG2YgJM4zpvsXY4Nq/CHZ
qrLP1wQPsMdpb63kMeQ1SqcIbQeWSIFzgunY2mweExviHVQc8jlFW8J1Z5PIBqkmHFTX50cxWEYA
gv1SumKfMuAnrGLWTRATXPb+7c0R6kqrk1al0yD0YpMGjf2RROxwEhj8qqkdEl0NcdttZPJoZtAZ
f5SaK11L2NBgjKVcliEk22hzd3DlcasXluKZgyeeCFc+lYVg9WOiTWNC9Mvj9xiPOjiV9o3XDxrk
jPmndIfjTOQiNaQHstMpRA9ETvSYzaBttAZO2JCY2UE/0G05NCDcigCtnSs+5O6QCmeJKJKnXMWe
SwMfK/zcqsunxV//l6ndXfdwwZx3pX/h2ezTE2E3DM/OzvmkrCfhp/hQCGFm1oXk5XX9G+oZVLIB
9M7/Kvv3PxxkUtT9TCYOwbYb5rB6YnVqRrcG/3+2z+tpvrxcHszzh1GBBVOoehRTFTXz6xc9eF2j
S6CVpBTa8SzN+Pi7tug89Jc46HJYjchg6cj5WhWG1DdmE++HNJhAfV2Xyyq2MeZIga9jyRSbeXLH
BEU2Vx9BF3nXuPVa4I8lxmm3CGiuKathvAibAdR2vNP5KaKS2h8Sz/AYbvqH5tLighG9sGGxZCTx
+vE4AeLnFPKwXclC8G+UKj+dhcpIHjs5lEPxPEJ1LgI65fWXtyBgzXXeQrKn16CKDxnT529ofbpb
S60FcQKmXRfQLggkMgS5eWcrvLRyEIcSVFqhbB688o14kjepnjAFlh5wSoXTKh02KGG07RZqfEtH
2o2LPNbmxfeamyBCjriEpZqNpflYlRgvUTX2FwZuOri05AqzcefZF+s1Fj2yOnwYUNcqeEbrIoDO
yiSnyLEoPtsXFWxJKQedrW2Su3hwzsE9ZwcEIuuib2ZKUse3AbuzovwwtOH4dfuUWljtPIaWxnlw
7ex1cFWTJGUDYJPAfDyUIRU4QSYB1E03J690+tnijK+ePE8hR/r9OlX1lx3qcJiF9pa+cA5VUwrT
ojv0YlEiiYV0r7hA1tLh97JeF43eT6Q4AfgC2yL58kq4ynvQmTtB3L5GYaq+EUdum0ufA+gEG4IL
bn5YsZmCJhhxR2YCFCe/L7bTgV6Iy+vVctY/smKNDNS9rzgTgkjWSD41QH8Rk2iNYthO2YDi97yo
LMFmZwM/ESOa1VIP1pdqKjRqyk14X+q7ywd2kXovwi17VyJtKZ8a+HhOLmAkiz7SoseyxwkeXs7k
leQfIE4o0U9Un7NGuOyn3JgcN/TtSY3eit4XUJM+7frJ6nMg4aKoDrehG2Hyr5w1gWxypDNBkdUn
fpzOubrP/K5FROu976gXRuVF2CjXu1tiLfABC2yz2ZIzgzEJT/lAorKOn1UiVCegN4oOv+YDidro
JNgTa1gF7Oexom+vaJYiY7inYTgRtnIQ4wv3KEjZa2Ogjt+vXAbUJudaGjVsJ6lEU2/EmC1GCuK6
6kKWOUEyCjjMJeqQhTL/USJ5ClzXQ3LlyzEhH1MsUljrVqK3HmO1qHDp4MrMVmcb4FpS80pj7tRf
BV+6x6ZhVhSLdaByOeB4CYIhYYABCPYvFuRxqN6RvyqLhv3sntkOWjAXrCZoSgBeMNd1OS5JuF2k
HRbQFn2v2Kj9V0vz7DMg7avD7NiO8oRkTIeJ9KIznO8U8ee3orhflmz/Ehg9SIk137RCwdAIGHK8
Ede9E+oiZuoCB91eJeY05kXztxXSlSQn+dcPEgAwSdcIi0XGGG/nB9jPDRFNKyci3erQ0JDnfi4r
+/zBzD6wUGQXVnbJaepw/q/ipOp7vqfdPzErTNCgbsbOT7+2HLDrhmHhhM2qifmzJn6SwHUu7pxh
2ec2ZOr1vAdROvuPgF5a0Lv0L8L7cbQbj/fjyQJ/oeKBnB2BN/VktaJ+DLkk/yFK38JiREPR5wJ+
BYfbxzz/95L7Tnyv6HBO3wUwhyS82K4gIr+Q0d26zEFyTY38AfpNmeKX+Qf+Dhou76MhkLMN9hZ3
XGNT/O4gcKIXaJZMOwIz3nOeK56oAbzsRWHf8TtldPFZrDuNDcMfou2AM+33e8tCKjnlI5LQ1rd4
4dFf1Ji54hP/5w+Vi/xQOTJXQZHSblhNVMNPUL4WxV6+zcECkztIcAHsoa2jYzQG8VEt0yx9IuXy
/uof4DddLhzSkX4gLlAAFcELRbo/IYlw3M+oi4XlQtBk5B8he3YyMwLHnSFNr6zoX8qX7VeU2ePb
av5St1FvWaVUC0wVxCyKW2qabCE7Ee9CvFsMB0Eu61JCTIYPLcGyyroGPe5wzWSGj8AQv96YoRS0
PCh3nwtLG3z2wUIEBKNcYDe/dZr0eUvQQO2NFsq1OlBF6k9CCKDvN6x2Rdts2z4iB3Cm3uyHNWr3
+2eVO9DEf+Cf7YCL2QY96Spd6+BLNL5IZp31hp5fh7D0vgHmIoRYcgFvb/n60+bK/eEmG2uFHPWu
4cMhoBYcHXDSNNFTP1buPx/Tf8bEVnRhLvEWKSU2ynzF/hj6sOabpujZ/Gw9t338U/gVsJV+fc7R
VUUb0hbbSc0bPAKusHVpsIBCspTVTYTpAzHiCih8/KPWTN0OjCMt57mZZsXv8efIHfbCfPXKqw0U
3BUmjCWVa5WG5WppGeNPXzDOuzxBXkYEAXAjG2LaGxFCE7/RMYy0WIru02tCe1XhvXgJ/rC0QKvq
zBLfbW37cNx93xndU/0arYjs5lM7OpyBlZRSLco0Ck3cx3hqx1u88xDo4K/UCf/K7Ohvtz47nwIa
tON/l5yG4jKxJM5bF2NHtFzOFPV9qlj19Un3pgeJckbM/IPZ5TnaEC5UpshaMEE+KVSJDyLUEV8a
i/uvpriZAjx0thmw/tkR6DpY0MS1fk01CNjqmwNFgXsPtF88rDSO08To31OKwKU+ENtLcuNYW2nF
+1VjHcDsUPRL8CN6ZPXoxbSf5c4ern7qzGFqCH5IcFQ5KYL5peQHvazhFnPMxhVV2fcLg6hzNdA5
1KQQINtnF8QgP9lX/u5//FsBtF/gWNaZ0NAax7ggM5Lm8tZWS7DPC9SAc52GbMq7beKnwJage8yP
n1JWowjLUXq0FQjghRQvwbKOPoIFnDUG2exc3EXdbx2XqTo7N2qAoobKkEIYlDnzVVB8f+hfkm9l
PPpiLrB1T381BvwJ6LLdYtD3CB4RgeV8Au83mgyCymqKJOJcsmfX5iyS0z4qnrBVcq8xDPZaC5ZR
fqxxHRsnHcGQ2/nI2+cIftH1egoTikApi7XhTNq+0XC6dIyj1qXEYhAGU4xVflY9QNysyaOce9MC
/Wgl72xcL3PYZ6alXiReEsKaa2ctK4fisZ0AvnGhNDVHYl1zt7N+vP4rZQ0EVZQOESvd3uaWV3EQ
23KdAAG2MIOUHAVwAL70OQ91oMTzUf2z8vGu24DWqoWrfJjbqrBMbX2fI6X34nJCIv7Ai4cnT1Pk
A2s3z7blkZu5b/Lz69DNngTKIvePTiGKi7L86GskZnzABuEU3ReeVa1PZtkPZvs1KG+g+4LDb4n6
75q+s/Yap4BPRgEgVyREoqvfQh6Rf93CoALc2Q2iPXDLdplI2KV7HBkrRwZoMMsnfaEmjAnaqEHT
WPPk7ISCc1vgzNKFETXUlsTfaOHdybqu3fdtspe2Ordj49RBO57yt9MM5ZKa/VsvZuQ3bt4nOClG
HprBuUI3LU0WqGQH+i0abKGDLWlTAwBgNb0DB/UVcL564raDiWgoRiHQoXWSFCLYPTQlGrKtXQjS
SopYvcSN4j61wkn4vuoDzMlLRToEXdDU6Ors2FGVjTtPo67k+nxv3YGoLyr4BxBhAvzpO7S9+Go3
1WEevxA4Xaz5LLCQBS0dxVwuxVKf89zxKmUKQG4+dL8wr/tgVG05zqKj7cR06F+Vn+0eeTW2c8b5
xeSaRNbYVj5HTW29RNMLAXIB3d0a/IbjVFCnrxRHZsfw9460tlzLsk/UFY7HPAmQ5xndRC781DSz
9Ks0yuIvQsFrQXrF9drTdMkX6AZPS+ln4ekmHpOtQ6IJMh6wKCOTgGBXipBGr37b/8dB0YDalJ/g
grCyWK8lLjbMQJU4ApgnRzZQLl31rUXfZAqHbJd5KQzy7mFHyMi3EuEOg6Hk0xoOQQ6hnbx1gu7D
W5L8D980zopU0U0lEJHNu7idLCfyOFaME6Eara/FmnhU6L4pwpSTDOYnKB0YT5sgGgGTVPwUFKO5
IHY+r1rhUHJUY9veJDwVeJbHeBUNana4qYUp8BpT5skbjYjRaBLpnnNWySPEmkWallWUMdwKdTJA
+SQufk41DxyuQ+jIorE77q3qZcBewIPyEn0ey6kO/rkfvUmQ8k+emx8RHv2/+ej7n6rzzRW03iin
j6ki1wT+Ml5yhmeQC3bCQGKPHBUkFqp5oW/qyXkGaUd9MKAUeI5qKQ7BUm6kD0llQZvb7yvJo0tY
Uz8JrdOr1Uc/ljcZyNlicl6KK8EsMdWXCIp0bRroftirdkho2F51anxbrrYI5kWCuTklnK/zvcBW
neE5PWhX4vuFIsaOtf26uzZgqAxkCBtvlNWnpr2HgtJ61B/PELgPuZ5LMrI2uWU83Sbdf1OBuTlg
Vd+vAzGNTltB0n0Ez/mggVvcK9FagCCIWVSnoixefcCRK8+jo/7zQr2hoyxST8le81hEEw3+VQDf
1epv/dCsAY+ak7Jk7fjEGiCl5Z6FTTciA4hXj0azN6NOKuCSHAz1O/pAF8tAT5+Ajxl5h9iMYLpJ
jot3cAUlKPzt172CUae9hs8ogW+NZB3kNKpifcVD7BDl76r84NSxTfOH76Y/zDi6+QfYp/ea2OoU
TKagGARO8Xlj+3C5LPeTxISwEMaxZJgVJg6G+KAZ1ATVuL6Gb11fHqXBGKMKoFfqcDU+8cYFXYJG
8+kq9rOoDEGnqk9LT6I6hg3cblv5sTmLbYQeUMrbtm4MjY9znFrzjtLta5g1okUNJVEEwDtCuqZj
pcY7kLo2pL2UnVMxaOqCMHU/0nMviy3mge7GHM59RO5zXAcNQD3m6B33tsMSHz3Ccf1ez3aGu2oI
yzG11mgsnXLaClz9ggqxhMKAS4weG3O3bX1UZCRurzZK72DEhuHGJdtDFArH/pA9TCfvimv6XIDQ
Em9ko/WRJKPmUGl/rg74G5DtSloKmRBACV08tIC81zt/5k7Q1Js+bL7KDgF7i+lIGGpvHU+Qmpws
7HbrYzsRIMbgWVB4Jk4EqGv91HuXtchqnUh5tCBRqB8DZYvn9XK9uO83lkS9H7MfVKHIvcmt5P74
E1QmtHlnLG5H4lSgZB8Cg5yic+L9zSPiBLue9brxeRcvyaeVXEiQXS3BX2RbrXsEeC81x4/22kzD
TVIkSvbQ/x02E0eVKBTN3R3EGAr0XVP84GLrsN3a8Jp/yMEEbHeBD/JdlkrujObmcDpnbVtYIRQt
iDq37VaC+a4IHh25qPZ9+hlLJsaGhUCauOOhyG++OJ9rJEcYM07n94VJNaWzEdwcVSJmjWOTavv5
6KMIf32zuscBgXNdTZApEKD48F7GovACLOmWoX4XLcJ7GpTe3LJflru78pwy1Q9U3Of91RR3dkhE
DKmiwNblfBnZQ7cgmvQZheUY0WF4bRjNBQQwW1HuTBln+WDzUSwl3hVCFG1nJoahm6qimybqFY7F
QYNss1b/cmpXiYQhLzL2lupeajNtP8aTL3If2aQ/1BsEYTQG/eXAiIigVA36vfJftxcjgLm6OZER
gAdMLrtgVU/6qY10YQnnAxH2hJ1apAKUtFAvXMX12Q57/f9dmqUr6KhsfNN+fGApvLdf5yW0BAct
RoX24Isp24h6j3VX8yntOwtCd4Q4uYbAWf2ob9WEsFL97N3JhNbg9uO119j5IpL2W6AgIq13J1sF
EF+W8pDSkzQwCaYUhcohQp3ftS1EKVKpBnpX/rUUO0pvvcFse2lpQlYqWLHvBHMOEzSC3lhuzfBx
scOHLkXy0TSLYMCJJhw7u9ni7o4H1pmGHpWYo7YrBAh86zM7lOTe/4o/g+mxVY3Oi6tvRyOs//Hb
xcVuU8TpkAQItDaVE0lddrmh9w5pzIDEyK9Tf0bw9gNzeEVhTmTLxVIkZ9wG3h0SywTEt1LZMdeX
NVKnLpvZKuY8Zb41hQJeqdHhpgBBH9KMlN2/JvKIBHW4mx7Ry4xo96e+UBTjVtjwnYH2ScqPFGlq
+wsUQzT0GKyyDAgNPvuFa8itO36nYCbNCDh80T5+5XDhS/UvNQR5lHvzkhvk8vturNva+VBVsdMw
wobdrhibjAhov8h5gOeFpC7CQdq9NLQvV9RnZcIpbCeEPw6IOs/j6S7uBpdWPJGi0kwPjwHNEiT0
w8INxWk1aTlGFFLGIfqGuVsGCPWASp0CLWJtl2rLCLfNgvZaA/AvWQMz+tgDt/THMc4vmk/UiZ5V
laDaPIcnnoRdNevSJ47FkSTjE80ju1Cl3cVhtI0uIAio/UZVzyBmOcrk1vySzp5kysV7QInp2Dtw
PaxPOaJrwVswYifGxzokPHA6BKLQvcTN9EIGZ1xfK9xhHJaR1jS17+1wij1kGBcHzmMdJL4Mz0Vb
8Oz//S8oOIk6HWoq8PeC0pBhYpWddutAKys5ZbQEzQrlJxSr5D3PPpZOeqjI2tdPZr1S0pz8HsWu
dHCj9bc2e++ZjZfAqmTUxxV65W+DW82rTolfmngbFJ7TGPgDNRcOb/GRVzRFnJz060d/LJ5aT4u8
xn0yDGw2OUMq5dv7Mb3+xGFeJSNzIzg7voqdx1A8l1t6ASRdgrJLyGP4d/h7Y5NbtcLyfyaMIDUj
77vL8NVs+ime9TuCDWWAq4bU6xBzvVZ6De8FnKMhUIU7GjMXzA0W0Kmbpky+kfM3OaHpk/FgesW+
NBPfffNhs/rGRaUI95eQaqQ79Q0CBTIIG3ARPax/jjQvZX1Qy6C757KVDdVWx5OG/QnBeJyMYW1x
99+wOOdicI7y+gG5fg3tSz6F2a+zVGnzWMw7y4VQuV7TDbM5T9gx6LvfwUt/kVLOS7/t4bDz2hJj
lshdy+dYPffj6BEWcXFqg7OH4wRKzvs/s0yox63FuzE21Q++p//kPTJjgKTJtnQ/5HagX/yFU4uZ
uU2JolZB6c8yPCdiTXr8B4SaM3V76Yn67yXnFcBELMTBITbMJb3AGdZeX5/0wis7Vkn7Fi5ikez1
DwTldjUNzuIHslwhLOg6j9BDNg6FjVSPLK5k+34ubHNblypGlN6D/3Ln47RAMlr7dEVpcGjAREfs
Gsacjc3XlOx8ItD8UI2PdHAXZs0BNt435aFNMbOjlwmIEqCZ9g8bFkhxkQ0Owx1iOAmpCIcPs9Q1
LNj9XU8PQTJWnN8sGJDPOBSR+P8fjGKBg5LXxt7oAai+vclmFMIsUkgl4Pdv5LD02ucAfxVOFiCX
wLr1aXXSm6+2MhUK3FAN5bmbVCaKl14Scd0Lml3cieGSZG0N4us6x3ywGrKKO+UGEdPT0Y+SVE+3
FHsrpqdYzspwME3kvUyBlm6WV3/3Z+2CpD+XKhBD+FSImpxLTaQQLhkB6NDvSChbq6DRXaBsWgHX
vb8s1akSFpMyndxQuLwGpzO2jXjowSKAcFrfJJiIOnWZtQpLG3MTmWBjgRUHJJDXhIQ11lOZnJgl
kbHIFha8vJtaxxmzNAFqUyBR4+j0f+ewtEAqR3mdLqwDSBtlp1ytQwuBFcrIdJ/u8mOl50j3QKZQ
UQMok6wvOCaXFYPTuMm2PYHAPqtMb8JaTT+bVwecFMY+rWYuaqdT6zDmp73iScsTFgjKXaiDV/2v
9a2qQQAulWvsvmdL1wbLnLGt4Tsb20DSPi2kbsInYI9P2S0hNJPwzcr+QL/1Ahswd449H0prmVJz
nHW7EAppB90saVGGx6nuwEoTrYE8Qq2Dbswqk3XdrxQISPqI1z1sWfk1utubaxda9pTmzvLLfCv5
GnyktKwQ1GoBGztWPIBxpcGfnDwf/l0qKwX3guEDxU/0sNQc52NaBSWLEZQ/Cx12E4uMEgGA7xA6
/QuyRduppPVafA4xv52d/mmcB1T7opq7QzkFfqgRASJ75W5DLQBC3OuocGpAdUMGdR6VmO1KNUnp
jA7hIbHHQ0YCU9/OR9HNADG76U88JmYK/cZFYUZrEbOQE5FSRNVUu+RIt3tlINJnZHdD2KXeSTG8
hQ0+s0zxuVj3gK6lcRibmTV/2PpinkaJ66oNEVN9JN0JTvI94IPM4lWO52h6MVF+tOrjWfV0yoMA
+Qy2mcpVmCjAGpuVL2dz0CAQjyVXd2ZOlhb8P1jnmLzHRhRtr5hTvwYZhoKVEvCbOZDz019ii5w6
WDiONHchyU/FbJaqqEcowjz97O1ApMw6/BB+Aaeos/+htULlW0utcpbsLKWKvlIveUEZ8fSTACPQ
oUEcKMpj8GkMSm/i+aAUMZvgPwXa63IdSoPa3it2kNqDgO5LbHuXaukllb8HDWrm4CyWvlcXL3iB
RJxvtTqdH+o1ka51LMRG0VYtHoVMTtDOIhY99NVuexMJZIRGvbULjAcPcqFuz3xwlfJBzVqjuGPR
k3HlrNPpe400jXMog913DS8SYq6Jk71Cs/IdCMpgeE8cWaWPYXuJtWF/R64tSoqtdcdZ3M1gByzJ
covFGJJQ8LTzqMtLy//fbFafzYsKZkSJvoN9b4CkeBlWV38YqwpXGmR4L2QwlsLkHDZSGNoFbnst
zoHNaR0eggz39PDQuve77D7p9iH6qJVxGMhu8inYq2drH+Sd3Jg/dNZ0q1xgSnt79s+DNdKZaFuI
cvN0nQyUuyipjEQQJ/TCVcSx3DYmYXzz0Afdf8idJtekbUP+zmw2ClKfzSVOJjIxJ8UOL5uXKGJG
uyzMMIXG+dGA9MJ4jQqu4UZ5oFNKby1qUHXGrh6ff0x8A5QW30xY4jGdHfGvFP4liSiTwe25qdJI
o0UhREKyrIH8lQqPPxNEjYCB+jACPdi7Y+rd/IGG2kL/ffb0vhUiesQGpiOIx7AZneh4n+/wNxRq
nehiC4a19QrosvAiT4GrfbeiJXCK8FkcnwKVL4rM5G0qyTqBMR8eMfxEUaoBZZCjvNUPiBzZO2uH
KibS3RTrRyN43r1OKTy19DKIu9YiWt1ZctL9CciNdvIWGiGxAZGVu9SFz797GkaHpcle/FCIokD9
vZYKRWmaj9pqTVxR9OzI87Nq38a1LYQSRBSDXRwRP9YH7uFGp/5OS9vk+/VEpLI6Uy1MmJTfWgEB
WuUsTG7+YzfgWcvVUw0DCtGTVWFUUdKVKIj6RLJsIsw7nNF7QrTJw0prlBtOv+h6W1dVtSAoSDXc
rJPyyqoM3/lLoHAcehywLOMra8WK1H4AbN7u+q00d5ES+q4lL5LoFzDkXqY8VlqMH8wGpHcssG4J
yi99yiIFw88qg07QCVnEA58Lr6z2jeepuz/NLkuf8gS+yxtpaVHrvpy+6rF9yQZfuFLUdQh63Upy
XlFJWExI54djUd+DhDcuTl41NuMATtEh0uendEBqANXY1u6R7WRciWTisCQp2JPrszxKY/CSroIB
+eVJEYlQNV0CUeJ9lz1fPU4nPA8NIaAGyrcsbTcdty95cnJN5+/qJgursXLUchIkw5RF4o2oLkPM
/T+2eMUILi8OqRbVw2FSzfw8vU3+uQPP3WB0m7sAxU1SXWxMLBpItQPF60K+Zmmw7ysWgIBVg+f/
XsQ6MFcQi+MSwJoTcANNqmNV5a59T9eJX2JwpcCzJpyFU+/ZMViobSB2poMYmBl+Eu5XBq0m7uOc
f8PSpMsMGGYSMj9pNhS3qTFfreiMqKMasIE8W3xYRyb43IPNQWi/+pYGJP8cBsm6IBleQsdqSyd0
JpOvEuj7juT5miy1Jmg0KWtVmcJimgXCRRfhVTXfaFIbu6YZRohbwVDEhq7KakcdgxiAzsI1nIRZ
STwnDH4PwkTJ6456UsTSdV8mhsLo/APXytfuzfgF/jH+rVxykIMXDixvGuU2oV1yZFCpsJOHVoAb
4mB9AiUtWHJZ6NnaR6xcp8IkMngOuXWrPSnyDlbsqb6+VeoB4H77yJL1GgpKDUZPCLhshKQfIzqf
CpIJ1UGIWlH+a3xjwf++cpzqvDeRFr7GAONerzyTKyFrLmugahruQJcOuGQHCDV5OuWUH8bxYMin
Ykelv8ya5RTDa+et9DI09Jp0qCBFeJjZK3I6SHKmCN67e3RYFp5Wwun7ik0CVrLFQLAAfHy3GkDH
IMT3GtHuYGM5JbgR1pcDMY+3ff9p3sZCFaVIuHTfULqPZvElBsLeQ+NH7P/0nF3OdANxHCcVnBxD
v6afHMmb5spYT8K0TxO6rYH6MNurDeSrXAQXNthEdGsnIQZRiaJnCD3S4ONuqp9tqKX6K6rGyIsq
xTzShtCzHk/WUtn7ehL5o/zyxtKgaehrnnCTZsdPQsqA2dqgZO+PjopE576bUA+bXCXcOVxNGRqJ
O9DUqctl5feVvQnlhC1GxXfxHhDGW4vVoHdb/y9y6jygvm4wV7jAqNUdpUgzffej8qJPEIHrTQpE
a32GHiNIC5rH5n7XLT15XW52VsNG24PHW4M5W2l+cuXdke5JYslbU9n+eY1rMzzTHUbUcQMS4TFb
R8pSJ2uwXmxgvNq00z3y+wuUzkeIM3g6eGVb5DHiVdwtCQbz0KWVFksg7r/R1vkZYw81fmEDmSRD
mDY+B2hPEeCnX7OGzgkjL0Anxk9b7sSUdCM3Mpgkkj/K84KR7/wKeJeqPoj4b81jDMOra+uYBK1D
LAFOzuZHEdtG9pAuJ0Dm7MnLltKU2+qSAs4htOQ0p/rQMSu5bKUb27CXHWApHKqex5ZTLskEWDW0
r1WG8D5X3bhH9CY9nnZNzBeUc08SbqMGJlsNjxlxb4pwMjcMGYHKr24/q2856i3nr4QQaxtGW/nV
nuX1MG561lab6CtHvZ88RtMq/sQNuzy/Anm8/kvQBWCFCzGWdtXVnjRJU5+WmYXa6ZFrhUGKDD4a
4J9RRc6Gg5yHsX5ejHOY1PH9SdXWJl6pUcgCeWNHYj63sx73gWO1Aw4o2GEkWvNG53M9e8NhzPOy
TKjBIZbgZCMYyFZ707F/jGkk99maaW9cjiowVt0N4eIkwPnYPIyZIuMBKr/tpOZIoQMriMCq4hgK
UhRQL33Wv7RaqZ+auK/xhJLmOh1gvIvRTe7WsKvfI+N+fwlDj6rYDvSPYIC36PkJrsfokNTSPYER
t4C/EtpV0PhtiKqdS7KmxouYdz7t7TW0AVHHPFt9F6vGouKRvqY/fVVxS29hgQmHVtWNk8VoyueK
ShaINXWjS7nqxUyQ3Y1Yl2NqfWZv4DKT3Drk+fLTG3octXRTujS/1rYTtLbiI+0t0Mn/hoWPEUMN
qK8Mzl6mjZiewvkapCcvDB9qlUfZjh0PyqrS4RGz73agqKy4DQQcIuIb54m6cGlh6YCzHVIwsEgL
TVc7NY8G7djWe/E7zSPfMqGvthYM7HLvtxQIylDIGrgL9sykiUmNNdG+/ZGOlBMuD7t6YrYFMiAm
CBdWhIKVsFQJyjAh6vqFXWjVqg1rJeCCvTNd/J1aWciBEgigtjw7H4bRODaBzjcSmi18IOKwKV5y
4ea+t5fiW1ao6Vml7cdMS+CLsLo+olnRL3TLi8HaDhve5MfQ0hTOQjctmg1mMdrvT1ZrzfbmI36r
cqVqFkWV87MHy0wCm3EVWYBzXYvR0IYQi8Ooeehre7cz+lm3YTYmyyikhKTmnW8iGiTBTTG11tPu
kgCLXZeoiYSAa2z/G43BlRTxwKyOB6UF5ZMHoOZqLL0ywerOlH0v+MIZfb2m9vtP2LCQHC9fFlcw
+fXSQGwMyYVqzr6C2Mrt05+jujNL134GfcO+RfDcUTEE81T8x+FzopAGthRkoorvjXM+jAcohy9k
9/juXYRVcjz3UGUOtEPSksJBtdq5p2VImqAWtVgWD/Ate/oxjAVFCMbUbyRDNtrP+2ojm2QRfSYZ
SQ/WynLTrikQx3qnfha26BLiuyK4HAPkRHvPzZ4QG3u/SHXmPYud7Xa9lq8Rscx8WzXjI5IF+DpW
y53pxgFCv+nomh1rs71rufsOvak55caocLoAFPP4kx+TSxYriupds8HNGJEUMFaI8/R2MRDQ0XOK
ctfNQ20MGP2aitVK29rp6eMqhVpB3EExW+UROT7fQaV50KNx5zgt7y+538COVG+MalYnjTZzTN0g
Ig5riID6kjBskpmlR1JsOqhMNU1pFIor1FL9glEqF4NlDKv1sIQR+HJKY/SDPFm8xxNmDmelrfRs
SLXm3C9+zv3sbTrFyh2ZmxCKXiyxMxJ0L2BiNP2pwNVjgVfEPwp07QY+sW003HnSpTwxFD3e+7D7
Vw0AYMfjJfEvTLGq0HZxTqHQn9Q7FsMyqFZJwxmS0x+5lv8FifnNrCIcqJn38WQxzpTo8YkCwLUg
rF7SfVWm3cmH8VO6bnILYLYnsSmwYQX6bs9CLa7c1jy6wnzm0LkkJ8vdcPoqsyKYgxGpnNiNDU1N
5xO829WiF7lGMnAYIl8Q6xbcSO9rOYhbxFX+itefTE+beg0DeuaGdVDz6DMT8MvNN/c3sJeGX04n
NN8OMZxvc9XzzMb5NshMp9bPdNPSZCT9C+NElbXPP/uyBz9a52RKS33igS1kixEHzK0DnM8WFxGn
9ViHYGyvlkMAAdN8gCCsJfld7P90LMMJgCSXl9vg6/7whQzocxBi5ooFaKr0Yhhothbhb3sjMtXp
yhHN+pk8sDMjLE3xy9yJg7xwg1yzKzf+GPG7eVLrPN6m7SB9YI5S7jnSAPSp3BZnJwUN+qWVYjBv
Et3htk8hesICg3TGUUDfOSX8gRrzLZOVsZC0hbOHkcoiA/Ekb4KNHGN5jk7J9aJn7zNpU6nvGzVD
lhMJbkND2+MpFZbEo1F701wG3O5EUCLcuJ8ZKR6zUwrobYpc6o2zm25fmOy3LNqICggk4TGHOC3N
FidB4zW/g2mAVWxL2kUeap2Gqq5j8GJtkprJ+x/g19zjJJfBiJIBV3VUrdcXHwBNVT8apIQbgr1h
LQprxUkKskNeEUQTfB2FtI+p1sN6GriXCX+nthtlRfMifzuWH5TVMqs+iRPNpIU82BH8AA7i63ls
fufIfT1pTSTRYFcMrzvhjHjqrIVGuqmjD2W2J7lLRjPuHuzYVNB9rHCiQDsgTIX1S1TQ9rEY/FGL
CJ6rMjHlmclRxtuSGl7JyVnGK2X+S3eL1eeYO1sxXTL1V6cgH8wwOhQStcFRM1Mc6lRRqhNfx2to
C+3OOkGbSkLmTa5aWgK4rvJXqfxRr7WkQ8qzNpzQE2r7It5exx3tWxZ1Nv062iQCpDVQNPU778Xb
iIhzg+kIdtz+boo8AdrgP+Uo4yOsuDpxAzfTkhsgn4mr/13riqV+5+M6TPsuZWcNgtrUR0hs+U9C
VaIufPJiQ9YQLYFZdvJF/CzY/0CQKaDndIV85c9GipOnrzG1L8CMDBnOE9cccAlqX/hmFProHTdV
WE2IbfXe3LSswISzxhO+7xwjuU0gvGTT2KGeCU53f/fguQGttXlqHC1uWpXc853zvehssVdi8tv5
7RDS0uMbDWYfsSJP+Tj+gojO9iodZ+5L0W+6Enfc8jRCrSSakmkApo80sHeIyPUUWpInLsu3aCuL
1T9RaxLK2yLoPJIyWyDaxD+v/yL6EiS310OSYyubz5arV4rWHJNtCPR7N/GCBRtWZGy6BMF5F3yZ
agCpU3JrN3dEtb5pzWrCbFNlMUyk7aqiLVjbvtZHXL3mQaW9Jh0sKzRnWlNBiBWMVGnk+LaUdF3J
WG3FxxTsNjLDY8I6LbLsb5bZPlLxgFZgzVVhILju31yvUneSMDeS4FVbIbsHFFastrhKLFeI/wY0
GLBZJNySB8BE9YlJXdGAfnpFmLEHyTozmRVRneqPdsRzDI8GSOm7Pgldbbi8sgZyFKCn0FqHfTEO
BKs80jW0fAc6AyJkMwS7DktCp/HSpIY5nCXMg6HGxrdNkYuM8Ft9L5hdais+nud+VgSdAUkMIwAd
+/mp/5pl0JWUc2ixzduJ3xKHLE8eVUm3QYmKT0kjq47L/Lmm5DBkCHr5dSCGZn1CTfddkDRrXkMj
7lXKLf3L0biL2rRVu3820zPnJlGgkHTOcufvNKUw4twj6mK93ATGZOzJ57wXk6OQWGjYpG03DkLs
HRPIlKp0JBnBktaHpUW8PSSQhL4q9zQEA2q3A5pqJdLolWDmFHvn7SSouTkAZtc4i3CIlzouhAEE
YcYhF+I+54eKJqvoqMLFx/IhNp0K12V8OgkG6+h64C6xpvDo670O5Z++imcNhYtCYLD0bzItSqOD
e3diolG1X38DYHQbbqmDFdqRaE0hZcNvHbESoCb66EqK+5AxkTQtYoSJU/0sVl2nM83M9ioITMbG
bjcmA1U+fOHZFVy2FXNeyJghGMJ1uFPNRdyNTdOmCJykpn9lRyUGvVEi5T6waFL1E6N0lkgkX9nj
p4aJaCEzPziZlGRMzKQoXLpLaxmgAISnvU4VaP4//FPhOQE2K/Giwd8ecUHAQbfDAN2PYpmNfvzd
ekI8EAp1Hbxh8UPuyohyIJMjaCuj6DBtqrjKD8T3F1YviqlfmZyMDmg8rcq60mwAeu/B418A8g2e
DA7LQDpnfebiuuxpzAesTsR+UrvhPEmaf9T8Ke/ZoWKLuXOHod5IoD5p71X5KRTHuTsgtGA8B5oX
sCGr7vaRRIqSbrKMAnJt0T1xNCpcbOgqT/gw2vK3v+um1a4SiMY+s087+jM/H68aSlV475ZAKb8s
BWOTlh9sXTL1bDDy+mnYP4F6L6A1NwQ9QYkOLWZgBv9xIvB+Jl5dbq7y+dCBI93/DC9gn9qrROCM
RIBuPoaxVyYfuDr9mnY/yBDWjrXkCmZrKv64Isrl/Km1qjn9vp41Teeljr/SxcdfO0HVXB4WjZ4+
loYr8TpwtoEMYqB6nxV9o6gI76CFq339dI5sbFQLvyaZj+SqhypSKO1aaIPVlBhnUcPdsdaYfMQR
/c3kLqRsU1xJv4Q3U68AuwIutCQQBL/0nBOkFSVeFA2IFm8izshb0AzngKlllBm7D588XpleSwuC
7QALzTYVpy91ECXDFzJBvpR+VPmVn9eiKBc9J2lEeS1a/d7oyi941tSNdqu5SYAZ1uLXhnVmQ41l
SCADGrc5niQqGvfFrkEAP67VHeS4X3E7YQhij3VBQVZFr47kGTTXFsh+iqCkRIAxCv0GcAAMiUgZ
toEsqKoWmGn7v8W+NOt8AQL5GfhmHW4ZMcCG1RQO4gsFCLCPADVJf/V5HC+nLW7gKGEk63HTytu/
rx06Z8lvXwZykSojgDPft2DmtR1dDdk2b8sKp2WXTQnux8CyVoZqGSI15B/sRUTa9qHvy28//xAQ
t5h5pcGCTbSKzosozG81olQGInkBcVWguxuCZB0i81QljAN8cRxOu9kkwqcRBUrif92Ew7oAXDAC
MJX5YphMjarQsxJa8M2f+Q+z296Dslhx+YU1E3A3o3aamymmL/tW6jtd8A36/7wa2JXaZFRMyp22
VLiNSh5liqU6A5nw+qPJuUfLbnU8j6VQ38T4SZxZt0s0jtU2lZ2lhffR0Nm8j7BBQ0RPdM0zSgpT
ySp+A6Y6o6u5e0PhQPrWFbrlJC4XbgYgrXeTwWC3ZCSuN4dUXn2GMZ3lwr5T4nAw7Y20ULVBRdnl
2W60x+veJ+uBRRcWUAUYrhwkRQWTLjl78yOobAc9MGajdNULZ16RTbQoH9LOin/yDXRXIprvGJFe
FcNaUmMS+LoSfSXTzzeOgSmZmqN7DP9iiCHFppsGnCeipLejN6DVcp5ST3V9TdlfJBqcSLfDdux7
Jg9riH17peYwYe380HifK/BKYr34yoKzi2HpV5ZGIrIev6TmqTCtzz7PhBDMfvrqv+zscNMUN9/r
sklONAzW2E4ovjIUfPbu3G0CsRwBwyTEahD3eel/6qaR/9X9ei1hWP30qCNKL4v+T0Gs69bh2GH5
r0isVKSbZMURITx0MyCDmwAGT2SYLLc02dB8Y94jsus+kv1WOWfYMRj6aT/R626pVytwFKTKWgX4
oTypDezQohoCvzAsWkYrf4OKyhCGTr+EXuvKsHYgEAbHfVNWyNfnPC3uipmebV04WVlVb5Szdep7
SW8J0v/9M5/CePq4J4RjejO45wDmVuFVVs+GaaTBsFwttz8YjHUIHPkqkWX15kjZLBdFe9DGI/5E
mFY8aXHoie7AYfehJKMKo9X6JzcocKC7uZtcg6sc7pmu+nXGxj7c4hW901qSOVjDqkzCMus8RtKO
TQT7sbF99xRM1Xv+MlV8y04GyhMVienrmyVGpD/C+nWkS428zdoxGM1s/LEeDYkBpgNmh6epCEDU
IeqsyHmJ9evvc+UaW84H6DMpEJJ717vCU7Tk4lr4ahjCZlltFLrSR58O8YrIjxGs1ZUKQ2/fBf2E
qIUGDEPIXJfQ9rdeNARL0K5xsOact1cDnqyK5fhMauN/lumKaF0psGwelWdGDh6VXLiKZkBbx0pa
j/T80cIuxar7JCeZ+ZdNi12OWWro7VTfPu5m7mZ1c0rfdLeXnjX0wemjE//rMxlGvM8aC36sNAjq
oR7AS89t2xwCiTSF/lHIKLJY3VuVdxX5ENKADiJAw56RuvOBIy23CTcYIbKQ3yBOaURs7CzAyB3y
rCK9LpWrdUkA0bTeKT6mPbxd+gzuAGRJN1X+oDVlx8sY9oe6Hks0nPyYDD8/qoFtlN267ADL7N8q
Deb8zGYqoLSaNAhRETBTBdwDpdjLs/pNhi64/W5E9LAt0VjyCMSByxvRpA58F2tinHj99js1wtaK
a4K/b1Z/XQggIjyTZUpfz8U/B52Dqe0/y4CFyGsPPfaLvZZh4sIMGXujGZCXajQpPv9SQY12pSQ7
6Yz8CF5+aCdOcrsylfZa+gAgzGex+pkHbJyPzvFy2FjgG/icISkpJNSSPePhHJ7cyo+efPejvRzZ
DWC3svhQVzEIu/I+zLYnkqRKBQLBURuWfZ33WdBQGED1Mb5928iZnsTIexXXxBiXAE7uWVPv/Diu
Jl4JW9goLgi0fB8TSPn9l+JrmQwWOkhmQ5X3w/n4d4QJfS/sWvpRR+AAshGsBorowGPu+dnIIVPZ
F9rL9R1LHL11Q6CRqni8IHby/PzwV2B6S9U2vabUFTYlvJjnvJbJIlha4dAHJ+Z6f1O2izUcPc6M
iSnVOZHTNOt4NatJKImqsVBoEWIPL+zqNk5pKwbWCdv9WSzBD08qT8DROXL+kIdRykf4oBiCGl1o
eLPNmWy7j6nWp+bsac9OENg+n7hq1IxIaIAriPHL0CKxAQmS1tLcVI8Fia0XHRheRKzbJ6wBtCgr
YkLjMY1TjHdfe4UTrQ8lVvny2pQ9Zysz880eOCnzYhW7bS9r4SAcHwMpcE/nNJKigP6qyxOABD0Z
nB/u5HC3pBX6MsfRrE6Kwki1Dq2+kag3j2Vaao0I6Alh8udGb993m8yScGo9EvsKCon5NGOXgPuW
H2I46jxPynoTWevA08q6YrSNzl8O/dkbjmUumKyfEmdEcCM9BJWnjRPWmVXUNszPKV7QFaubIXCF
5SCIG0NHf9KnKefNQo+77e90vogEm7lUnZXZcAquJSki/jqK6H2jynkM/Xq/arCHFaNBiLGNkwxj
1oPOPfVjL1kONNwfnXiz4q2ZvIJXVuH1Yl9QMDxWhghDtrs19uMDyyhZ/wCsMDpz3xciHto3bbCa
AM5vnqyLrhDLndVWcDCFw8ck8PuR2uw2gF3eEcQGwz3Wid4buNsn7k2hVDinUJ1sjWihN5IfRcLT
2Z7LXq5H0YkXhYTVZdK1Fc0T4x2uWN3jDAxoZw0CnbSCb9ryuUB2Ujrznf2cWfIAQRxcxDcdto8w
VvYxs1k5Hi2E6+xmXK1uV3yQqCSgCsSK9z3BSJv+wPPflpt8eAal1ec7ZTLl6VgIIWCH0hh5/EYV
g9eKY8EMQctiAsn2osSB+2ufsl80FLZvYp2yO+AqLZOgzBZUYrKg0Wo06VkByM1uVY1imjf9rlKB
+qB0Xip37Z6GlHrXxE4aX5aHx32iB1rZVLrZvYjPriKCLu/84GKxcxd7qkxpUtAH3gUiTNDkvgFX
FOiWLfWCw0r2Nhe5iXkKCaJ1vRJaopTZgitNLg0FmnBI387cb1UGUQd2SrZLv8p/qCYWnCFb3ghM
jfdVZhOkpiRxvbp9tEJC9jFX/XSnu2y9GAJt8j1KEh953fkHpLOibBxhDZ/Y+Hl3By4yA7RrNDXA
GBDlhgrMtAb2Z+4sbqQsvB2Mg98+ofGlOsA1gygmzNGXAhWUm2xwkV3IpCFFtSUVNrXaKXbddixI
ptxJJ929RLiKAZg83AQVuzxuKS4IjBdNvL1ZQxGXjBhtwCAINAPyW1uFGrkfmc5wLW3/EU5r076R
WO3kKi/f2nikkTb2Zu+fdRNkOM8uK8rHq+d5pPqQrilp4INTLD8TRVcpDUYy+v79M7oFlQIxy8o7
j8RknVfS+q7aLrfKlEKiqnclCYUoqXVeLKl7xFAVQtAbqxrG+RMdBAq14+u8itpHF82IQ0QqPQk2
TKNJdudUUypmc1RdJ04B1c9/kT4TQW5Pr3yu7Yx8iVWBQdX9MQrzYT+5d87OqshJZbNM21/ZtKjh
eGwDJ6UAmBfP32rsJquuS5MtrcVbpJ83EVhcOBiwZmi2thzhb3Ki26Q1slJdr5xrN0w4wJkPXgxm
+uPJHbZa1/Do13C7gkA/ThesATF0oZNC1BgC7OCoTh2XICj/BQBPvBKHpnKw3YFpWJyawSrzflnZ
J3G2QuYN32CoZJJ+mOR67G3ySo/Mz5A5eyBr84UMQsgta4VIuKcJuNW5Dgr9/UeQTor99bt/o+U4
xSJsv2nkBYqzV+zzUkrNhsWd4woDyJRebLwy7iHndmKz1C5SaB+S/jhpWD2WS3RTHdvrhOJns1sm
Uk6ide3ivPdApIKiSKNCY24VoU3Un42DEl1G7dH+STlYZlTHB3cO3aIqjLwhRb2csTX4MTltmqho
qFnFwRlMJgHOsfiXIdCiCpsF59GeaqHf4We+FgsNz1DmXuJ4tih91TVJ/QgvFOA2nOIWK0CmKyHS
NoFHqXrUBxSa+mRxYgxdmXauKb7nyq6S3CEkJi10JbyB7s7QSPEfnOmKqacBxVOKxfgH/e25wF0x
xgJkspN+Smpd6F2Eqr0MFwYJEoL2v7SZP5TOgH9JIrhWhTR2IoXT52BLLVRRXNy7eCty9/tIO+kN
aX3GVJA8DnTHxnYMSwm7qKQA3lKlFlnSX/VPvaTLJybbsAIOnTkwK3Ft/6CkCpAWwAQ0gtds+HNQ
qwyv9Tv2FtEdTxgDTGGaKg8lUeGevjoK3R+6I+ohukZ6gpX3zZpabzeCfwWRxUOUiaizP8WVisgY
HoNjFsg/Rhl09O4cdPYNtbnuWEcUYKbR8bED9eHsQMT1sDPLDxfD0z0pL3LrYH7jgF+rPzggnmtg
IxE8/AuKZC2G/ia/6QJefJN8CwGLMxHSYQL2NG1toV1Icvm3dM9RLq+8R052jkpHS6wJ74DnEMox
mVr6ZmJjtCoAI/dayngIHOO66+3nAvIPugn770VaBMPCAbQNMEdw1WUknr6CdaEdruJprxegJRA6
8Pxba5EZrnLOG0bnq3ECfF65QRccY7dojWF2BS1gL4eUsLG8jr+CBTuvzgJd++xDjYThmRu3E/s9
1gHpRi9Ihe9GBFfXwRsWXs5n1lhBdrzDI+cR5lsZhkfhyvcfhluePH1cH60fZJf0na7PWsvb/Ju+
/9G6ZJUgQ8JzP8Zcra4RiAOzgAVOU47pfrr4oPkqpUdGQbeyDM3yfu4cvjP2Za9kKDLFOkzsvI1C
vRuLo88tY+tm6pkmw1yEztchN6+Tko+m7hL4ww8p0yjL7prVBttZ5eJKxiHHkIsaRcWgXMfLJB10
bcx2jau+dFlnbmGiIEEUuOneNh1EaP1liAlpOYJ06RC1Di8cntKNMhtp6I8C6ZGZtiPgAyoiQtLe
y1zk/rHrTaGk2ulOEpRAAcaNRQ21H/bqllPiOHScR4ktZ0uE1owA4LVgtdjYuEYfP+1qefxoRqGV
nuBCQBtxq5BqgvZxYFL4xKAR/Q63FQBq4D8Qg0T+xNev/XJrC6vO8N9vT31vrgCaQrUSM0PszyVh
Lu6YxDWP1/nAVlJX5IzhSTiSPvG+cWTvC84B9rnZZZy8AASsR2t8jHu3MiO4FWP20divrGlrlVc3
JZOaJqhpeUYgyWMOlKvv7LE60xKxgURcdoIFdNP3tjtCoz1o9g2XSfuOxe545iBgOcWPYYR7/8Hf
KRqIxNUn+//ylwkBtXLPGaCn2dZRQYd63+lr9zLwu8vc44oh1p5kYA7s9dcGSHcmgHU8MOQUC6KX
b+oNzodrvaYjxv1Oqc9rvPrJwhKJKhwLklBrmLqgWEHVJ4vI6BFb/3TB2d3fAiUI8L6ncYN7Xz2N
hpcCf95N5TOwtN4lo7EU1NrhlnTHU/5DeNAK4bLZ1gngLEDk5a2dWwuFaHDHQSa6aicCtyJUeZgJ
2BdwHne14jB+hImXbaUxr2cz7XFqEkdWV1Wx9EG9Lu+Fwnuzho32RpDNYRSR7NF/kHCnp3CGmKPu
C3k9diosXzogI0b+toJ7DsEt5TTgz1Yjg7wwcHXigAl9xh0DLf+sZIxmVdLchA93mv1HTfQLLsKH
07JyZyfepW1iYBiprHcZOqjQgtYjk/AOtixQ38StQmIqfDXUo5NamrZp4V4c/mxjEgtQtcQkopN7
m3eBUXZp5YgxERW2PrIpkYGX8r9yPWnkf1nggkroZGmnY1ecNZZKYOa+k+RZ2mbT+nQ4tGpx6Zk0
U+sQ8nJv59pAOB8EbjQjsznW+4wtyxKm28rfzkerChVclGVDDymW5rHZ328gDgx6u/SDyQ+busnF
mMudLshxrsYZC0WjilBb/uOf1uawhe7foPY615zlajaJItZz3ga3mC44DzMfwlY3AxOnyPoiS4nS
EYxpmsP7ytpn15zMJiEZyUItV8zfooA5OsLCN9xNn3EgJVPM1ff4gNHKVxRGIrV+N1pproEvvWfr
HdBaKrKQU7boz+lkbEdUF7a4FMP9nX8yWYlTVrk7zLZPCvNVKAIH1viEwTuPmlcLZXdknEGhr3vE
TKIu+bMnw4hX9rEQT6b/YwCcajZ26aXuDs946aok23CjfJkBQ5fKA0IdKGCSvjbIEE41mGDUuHwa
iz7gKd5lQ4+IyJAgvLdRqCEaLmla3RwRJC3zRC3IUF4+j8WsP5qGsLmzHNy8YYc3SUtd+B9/HmxN
hdzG4LjoY6ytEHHQ7Ipgs+OHkRNcBN9gLzeJ2VsKktiXWVDm5thw3nJ77fPMc0w6a+Z81YU+nN+I
3KMypoM5F+2lvXyfZbakM3Qted+4h8Fn0OmRzBx6ZaQyJ/ZwuVZ7/tKXh6jI23TzgIOKobKJYrEe
WCl0mNVBb27IAeKvw5cr8CC59WfsQeBNDztHZ/cCE8ygWPSyoLuU0FWOnJwjm+94y+0GfZsCmi0Y
GQD5ydged/SXeSiYL1u9WVyhwelzBfLZxw72ELQqNe446JJ9yIKq/5KXnIXRS9pZYE/AYcWW0Fp+
9V/IiSWA/aYES2yp0rPHefFMfV75NZNAMrPzj9moXGz5o94J7oCcMqFWEYUBtWDEIqcqns6d0afk
YxV3RAR5eWCPn7AU/17OdbBk3ErMam57FgF9LX3Vy2xJ4LZHuPP7NGFJKFowfm3/OxBNSHOXWd99
Wa3tvHdnLz8lMpHKSrpIcDZuuFV0maZWzEdMc0BegNv39vNz9nMlyv35ZDAqon9/lBj2Si4Qlmz2
qo7EazbKPLGDguYA9bZWYPiPFXhgpialfpvYq9D+26kCdHZvOhQ+IZSSmKRfbdLR9nQeM/TChy7p
3bUeTv0mgkpNx5gqkgltxuW1NIYbaJBq6ImCFntcwgbsfznR6/+J62BHiEOAtlnj4yjcxtqBMjd1
uIxfK2gPINz9AncR9KNALBwrAfNICTXlP9eg8dmQMULWCO93coKJ9Ks3YvhSDbVwbOvgYpDenrWd
VNy5HsypPKZlCacF9rN2D+Cz7NCda2+SZA5N/GRXO03AEeMALdFFs0GDmtNTCWLI6ZTU5eY/06nu
000BSORAnwmKKkM9tx3uqhuJncf8Uiz56Cl0K140g1wj5V0mYx2kSLmcTBHTs7xgrM+mbKaCxo6z
frf7B5WF28sB6Nr3VUe7Jlh9TvQb/eQMVnKPeh2J3Dnv4tjXx0ojbK23ZEQddG8LxE324k1tynru
kP4YHwfs8eYwaIhIgQPcSy3sb1Sz2SGYpIGQ59cxOalSuqgWx55WGsvOLUsd19VTRCj37UrYWpp9
v3oaViLLEGfrhF+AnT50XQtqwjTJuoVV1SNg3hTFckYqJnFvWRDqHyY+tYGqAOQpCXXkr9tVLo7b
t++qMoeDk7OtNjOTwp674ZtpCAKcTjhXdtOrct82W72bwXgeycLF0zLpQUH+MbS/rlAQWJ54Rd/R
J2UKj7fUH8x+aU5jqP1ZG8QcArGih+OpkQikUTN40un3KQdDyprUUauBosuYLllqFqz+dXNSq9cp
xs/OWeNgPs//+wyb/AKOU+xrs2dolcep+oqF5PrJCb51a9e2vVQ9vv3Mq8Hx9EjM8IJ73iUnVF9r
wgW8vaDM5wNaueGMj7/JqImQjl2icURiLsFtBbRmgoXiHWeA2DPTRUREftM/5fnpMmCqZbJ8ujSi
XxPNSaetMpBVFRpDYjcwWyBH/RZJI9Iv8C0/rYgDASsG9c5L19KcixHEsExqks18EjXEyAlwH6A5
OCpNMnZXjj0Adv12l+gENDUiY77gD6jB+PhJKI8ItRvsRfVPfn1Nlbe6XsdDkunDN3gx0NL06O7Z
aOZH5LVZYbBii4PIth2T9IDOZfQQeVAagbvMpSyhRHCFe1kRLo7AamCpWjlKDrY+eDNjKO+y3fEn
XsI+VwNsXdsBURyMc1nUOjxuZ6AvWamUCeN3BLd3tCTKen/+UFs4yeIRuD1cwoRC3bhcAwIloMf0
Gvtj4mpw6Ubk5dC1pp8RJSKsMBnXlCN3UyXLLxj3+hoW33jNeEFyA3CzxB5WCOhH5BWyQeGte39S
GPNvTphrj3kBHvrQ11XUYew6XaglAhO3HKH0wS0TdHiN+hdU5TgEiyAutAwmfGU30es0eY+rtWmG
YUcUyyUaMEgTgSVFQZoLcpOYYpI7Jh449+viQ4+fEwma+UyRVP2QovkqPUNsKEvguz4E/xYlC82B
da1tiVgvA4TnsGbNRyOuweu58U7xdlrHL/KffCRYSv8kXB7mx4e+NCy0vh4pBRNtLD5HTZbY0P84
gHJrGAH/36rUqoCI43FqP0dAsFLM78MMecf9/lwQKZj0Yu16yGWlS/oeNaKGJBWWSe6MOj+7SJ3d
kzlB0GSvpNvc1Dde6LjDEEa8bS3W7RabQGR+9/80vAJfK77jaQusmtkXVy7QkNZbDxz80kOGS7m0
ffhgPz9A7GQYwLP03mmSUzVn3x5Psnmf0B7RWd1qmDdVkZwgCwXW7brpb2GpM6B8L2a6wnsvDd+8
R6l2VXD8zCTvCrOrfubPHGzT6TOMaxUS7GxTMQDJ0Mc4KarlLG+WaOEDx3ZPJ9ihSSnFcAS0y5q/
bUDEwSNeBE+HLuHGLhRCfMbXugf7iWamO4Y8kxSeV3wfli9ajqRSFF5J3koWXOOqdfSaWf3Z+AuF
cEgHv+MDOgY1FiQf4pp7E3pmPVt90PBXYzF+WFDTDmrS/aF8zlidJflpVrLvq2qMdg/zwc1CQI/D
ptRBLxRYUnFLRA95larEdyBV6oWgNMnTsKwZ/5ra/zEzyr4pMsBq/jtuCWmTjOABIR14Be0ch3JJ
9aaZBTPZxPtnm1cFc2egjGjs6ZnfWqZ4odFNKjQedXmfbj3Z6fwDARUKdo/ctJk79REhJhD3u8qv
9CU05MAA+TScWY+7LoteVgvy/j3BQs1mu7UPkDD7gVWar1tGfiUsX4ceAou95O/sgW4rEtV4548j
HBrxU/Lkl6DcwQxqSSTpEbNbN+DiyQsrZ7zHWookBd/JDZy26gLpFpfG9K2efgrPiaZFJjTAHL+4
FOPpYNeTP9EZ2wlJVhQiKRL1tBpN4XS3BTL2WtqVCtE0T5I0jZbtQdioYONe+JOn1rMvh7dwLMSL
+GyQ9FwA34ecXrzIg8LvOhAGVZlRL7M7cc9L+chBKm2UHxppN75LLdFPBuiULSaPivvnQz1QYdO2
hpZjhHaygCJZHV4CwwXK3+imTSH5quHasNIDu77HBQN4Re3Ocz+1lBmd5HDcq/etLp2T61cQZ/sq
kHf8bcK4HiRKWFs0fhY7O+emB3RSdVEa1G3bbkjmbYiZcIV/eo6ws/mIzAjt1w7YVFi/DRhImswg
+9u2ze5haKJMPwWXZYkKof+Di/R3MYSqNIa1a+w67dB7tGROYtL7hOLugNAgDuJ0ZzGSbPJV/TX+
5MiKjdsHo7DSRE9sD+XLbWVY/UQI23zrR6gkijdskYD97BzvaI6T9KYB41fMiC6N3u+5a/UZzTJa
6eC4qD2EF8WRAAjQ/xPpwYQEjHhjW7V2LY9y+o0Kou5nnIC9LX8iDVWmQFF8wm//DU/F2zIAYCjF
6/78ittYge+4qPheNDGvcLq3XaJxxZMDxCTTYraVzzFPOoQvga1zfi6gZNNB9VYE+yeTd4+rv27Q
vT1V1c7a6peCB5yb1M7gXZBjSIuRst2Fz3TPEUKz4eemL8UEVwAsh63cLErSBch/oPERKv8OI9A+
HAp1auc938wAl7cwYmq7hDUhBZrYhGVpxuc6L8pJWzr52PXSQthXk3ItxAomAdTG+j7NJGwj2VFr
UlqAHxsMpj9b5dSKMU79W/hG/3L8qQKbTcq6CHG06E8bk1i4ot473hH737lHkB2NCRcM3BJXgQQz
FjoeTo6Skt5+KF2PcEZjSASmT73TnSxBh4njBBwpAJhlsmOudTWlI3BetBCfdWJovdX720Z8AACw
Qh3SdGExVOxah1qYY7K9MtiahCF7FAmCHC3+j/qHOj67onGm6IUcRQoruTFqgJ0Ow85yramWyHc9
5Ui1ZMqqUsmhzB7NTEHkakfTWNUVhV078qpOSBLWopLkjdAO9CH0MBs4zEB+pQpy9qYag+S0FXhb
XZBPRtuuKaSl2M5157sbkbxhdL6LMRBzf5mtgptyvVoKvpfj4sdZsbKYrflfJVWhXzAVR/Jw9CT4
b9NzO89QUoGw2+J33Yubdr9sXlkhEcQTHJv/0MauOBex9OjQL1CIyrgldq3LRvaSQSNU9FTBOD0B
HxTs9Cl3XdVYxHMweG5yEKruf+Z2I9W8Z+bHjRwko6auvYSD0XuQavsUMBjbzzVQcRuadH/H3F7k
vnYLCgdk3bpbvfCGiOYJmqMDTnu/25Hn/qYJV7szQwz8eFk5RoNtVxCFjnSOev+uZVRE+ivhmtd7
3tmbo0+Hs0sxRkNSbrtx6V26OOYWaYWphhqQ+xGol7yBfjUY2mVe414Kq+s1PzmjsCVkMjBiG888
hr6f7nfGkdKYdoEMOVzhZGHhcevIW9AKZTiNMeemNHVKoK1TLB/YBVJej1farRTTy9H7Bj+rKRP7
47ErMpH+VFJfkCa+vTf8NENvIbSWLVnOlefhEplKZuf0YFM9YUjC8CcLR3tfnDvqDxXgKKgoMP+m
QjRtrlbi3fAMk1JbjIN+TZyr88gYEUqqlskYE1W1/k57gY2IciGUj4lwUKkZbizTBH9BGJlgtRrl
MgimONAfdrshNgjPx68fTU275bmxAVK+SI0s5/vmideV+jbSfCoJ6benE3ull0gqxNjyPeIJAzXf
lhB3NBSqleCDE7zNzNlt2dxzoZtxt2mIGNWYl/csRFy4ka1amDlRbMQYwFuvDKQtXxdEKT2VM8qh
mqjZ26PKS+uUIsQU+zWwhygwmBHeElSXaPp+mAev6g/QiCjxuRPflbs826aXn5+I2BL4w9Wq78fz
ina66Jv4dkgBjjq8uBBqAPwUjps5MiLRvEDaO/jVhH555bDEYC2K5j0zZD07kVwnrSnI2fCAZ/XB
GWoSeMbkXek3xZTikbL/le2yXNHm+UzekEHS9yi/TIi0AgB7dH97ut/mkkk0eNykqNUxMzyeqlsi
xkAxW4jpm5PoKK6Y3kvhfeX0SwnSLZP6NwZweTJxtlPnJi+FXff9S/6BJEMtHOLf2bZlk0uruxiz
3pIj25EWhKr4LKqm52BuY7unAZVrZqsMwQ20gUJuTde4bW0ifu5vMiLtDQeuk19aCauoM5DrV0aB
pV61Ybix2uIamplj8pFDcFyYmgTgzkpdWo7O4tz1t4xfu0C9ve1RV9Mm5HmCBquhVka1p4EfilLU
FyAsaZh+C3UmH3t4euoCOBmUAkZjI9RiPSqaAhNq+oAIjcFiTRDhpSQWQX9rtzJ6MYGaYq7lhiJX
K9U1uTiTPT+4RgLUnswArerOwUlehkghVDMD9JpGlYJWx4B1lp+Xmxoi1zYR62t8BvLT9gWMdpFb
3QAElJuE1M1DSXcU72Ro5VtY4YOhkLIQbtXy4r3NJjwTHOMeGRo3bk2oHUFqBfaoNMKqE5MyKkZG
HTcywUhza+83Ubi+2yYG/uuu49aM1jwh6fn6r/XahRUHNLd2pBkgJT982FSYe/GILLeX1TxJxK2k
v7LVn5yTCHwOwlHErWfG4JjbHpsDi1Qf9XrE/aTFN8PHAxG3tbV59WUQoc3IA6zcI+wVb3/WjXrB
uFK0oA8yqRJEYOJVI5CZL1xdGgV1LfG79fGJjFKs4SbrD6tUFzICMw7K8zOn/XfhML6ZuQn6Tk8u
4zfdik43VrCQE5+QwycZTdeA4KpNskhNHaI3jwkRQMLCkEDB9o4afyMIzRVJzHeqSPHTaj4EKdtW
DpAxfuO3GvyREG8+R9wtlBIpqBVvay2chtEMGYrKVLwZ1u58dkoCoXDXzBRbjVLoMXQJkV9frwUl
dsqr2Mfwm9N+4R/+QVHckLZ+gLThAx1wAO2UT0sASxOi/jZ5CEob2yfoVyaEEgAKbzRzzslx5SV5
54xgzR7/m29ZWPw6y7/6hkZId71GicfkvOHF+wwsPdHjsiscRnXDAEklFkJfPi9lIV2+yFf14MI2
OtAAQMyoJdAjNGWUT+rK6y1G072ToNdhRr8MWVQVBV7w9wBe9hSGtYmI922MwB+mzTtSU8SR3dgX
qW8Dw4202IMdkLg3Xt3wvktKNxzQMf5lggkj5R4IldWRLEeUusRVtT0wc6s385eJ76Gk7Z3bNTDz
jj03N4EBOwzlwIfY1hRVrkOZKke4XxYcffIO6TW7ODIn++xF2TXsIGDMKPMmRFheRV0tg+PAJmwL
KGsqN2YAEkJR6gOS6/eRubK0fpzM5TSMHmdT0dACzVgJob140od0YfeqYqG1XGu4hgWILkEsBc//
A5Afs0gvI6sZ6o2rB/ykX/Q6LcjAkj+a0GP2chx7wL9VmxKnwRIWnSm6D5MSp1vsJQ/rhcl2SXTA
1sFpT5ALq4r9o+bPO+cDzjqvn+Wxh1IOYpKpSfI9P/+TN3q4OWLzoaD1SEEwLxLk+QKCjC3hMwUl
d+JHWJlulA6VM6OIwIPMqTHiJp1p7t2FNZUasObMRXssa0p9HpRKlIWe5CrowszzIVbzKv8ZThFq
blfrQPZYmVzd2PztVWyAQ622VeGseC0W4PWamvJ5t1lKpBtBtQp9mf0nzVSCbjdrGxaKegphpQoT
ZvihRKd2N+lxcpF4asay2PyD71YohvXu8h6QHpTG/fHrSt+OHA/TeLcI/Ss53PU/WZPeG1gYSysb
wcKwHi1Hc9gy1egEZv00tYBW+qzpUIs5Xdtg48C4nwsoXisHIJNuNikC/uj2uK9Wg/jdGQKeMCnI
KrPitmWvIn9lrx6C2YzPZqhb+H++MHSYCf2d9H9VNSCAH30viUdIlcivz0S8clL+uGVPoC7aUo5e
hfbMoP/MoqEnUlo9Gp+9YMbg2DhcLJgsp6wElwXNQWggqDw9MLhQocrqM11RYv72VYZwflYaBUJ1
LG5adPVnhMZUf0lKSoTLSs9tn8N8Zy4IKl7pNsOloSW5lfB3BK2WsDr5vaQN0YqVbMPT205sZ4SR
zfVxkHpIu0q0akhApSvrGgWzSIckznsYbAUFsBVJ8BkECtbJBD5b98nUICG0V/Y+S4byCoa64sG2
ZIEX/EYGnj4VjrON3Ghq6b8fqunBvbXS/HAUFHGQeRwV6NRy387K0ZndX8ajThYLb32JYLhzyQfC
gvnJBwN+ZTfG9QsN4op83EikbFyabb+U3y/l8MVf8ndRGtd2qwwwFLvy73rpvsvGML9jxGf/G/rj
QziRgcGOV6CbiFEx+3nrrzDxQix8uEpaOyMefWLRVN+Y4aLOOlssBIxcTI4QKuWG5vjGHolUMRwj
p8bC5CDk052vozK1An3w5915djIkRVxqeN10l5uv68jUrb28nz7yQjg1yKSQuMVziVzVNyX6u4rD
aHt66OoCCDghhp+LuXKP4gb7wC8wKlliH6UOn92Jg1B/CtbZahUZ4m5sHR30TrSx061OhRUkKztO
0abPov0k2+EJLJP5b7Me6v12VYxwB9AYOo7A9JOj0dFvj6YkzrU4mbHVYp0v4/s/HBrob9/KxU+v
z61jSALGNff7jfh6NY6W2e6BHfB/2ScxFsJ0ovUsBwDFKxQ5HtXfzL7mGOvuRPAGY7KzhBZLNuDo
DYagJuzyaZW3+fd2eajIKPf72ZGJrmomyLNeP+dXb6DJWI698t/giB2XQAjOcTnCIiq/yxNyzLTC
fBIokHqxAdSV+7JQ/s8g7/3EwkrTzVFWonmOQVZt1sR9gc2s9t3FjdpcAZ4y1ojFcwVtQzfB31Si
HzfTOJSeA9znPMwGgKod5dyYO7kJKO42DSA/+8urNlC7lRgCnDz3rSizGC3Y7FeReoqdStnS3vU3
gF7oRELpDvQj4ponUdN5uSrhu/BM6ZSAiemThOAjvJAjkZe5ptjGHEMnD+tYti/z1COOrTRfk8sg
aaVwyHzaUVatTuDsAtEX7EEPfeC/gynl4tOi0Lo8A7DyfZqvOGTD5DA7Olxkv9/z7m9kzDvFrr5S
hwzxmesTwDohwb7gmZyBRAbe7eyhb4Xw7q+QIeTQUAgqF9qVqKIxVZsFDjpvL4ErBlhrnhM7HX/j
msTUr+zijxK35u1AVjLzKMMQtsLiS3XcG+wYqsun/5a88bngEQQ4xU4Sv4oeLW8tnpv7OJYdmOMJ
4aJGfDXfsYE1+4Ycd5NP4XWVv19Y2kM9A3dDjrAw2+zOi0gEL1rMHadwk0Ovy3gzSSCqV211/7D9
iw4MjzGei4F/qsI0tEmd4/SUDVlSIkollvuoXEouuZ3M4rpe6bzChpOYWTwe6qexwaY04UFDYzTf
BDuJpnPAy9Q2kTh5KepgI7eaSaszt/6wwEdiFtCdPWtXvcsil5elHpPAjjf/WMh5vEGeHGDHfkVA
TX8ZJ7hz1hKGD4rGu3GTY8uAM2DI1E0NMT5HEuqJ1mv2dZb3Ezs1RugeENIeUE04clw/Ar5P62/r
Y0hCoI7Jl7agrZgJ2SEqAl+MzJMv8X4JBfk8TJIAVbesohFsfOJlUGqCXEVlIFyiOs71ywFOJdod
jaVHheXiqlGnjyOVbRRKJF3ro+Jksm9pVlH/yUhGnNyM7iJtpz0LUD3w2WF3GpW4LiSO2BEUlQ6Y
A4oMKvfQAG6Ej5rqLNG0fMkWL2uC9+Qu8aruZw03wN8RZNQwn2hUkVlesc9PRztPe/ePJzGos+5C
bYfOWM92of5e4DIjvOIYBfqcknGuvm/71qnV/XW73w5zAyemsSHy+ZZ5FFVmZClOPAb7CFSLJlvP
rMx6vEGJbTSw4YzN5XvMqiyjGk/YqaSuRVCQKB1bu1668qxZwujGtlLl99UGWsSDnGydJgRa+uwE
Qc4l0iQglrnH9PGc62FmAOTBeu0+p/3C0YKALfxlQYlJ5dfDuzhHOEyVqoNL8HqAVMU4irnKmaQP
dEMynpGpIFWWNx3tZuW1C5TNYapPPibycKD1cBQkGTK9YimMJqvxbgyF83fmfuJF4KC0xP9H7Srx
JnPrMrjMCI6OeJyNzs3INx2x34+IrIXlBqyRuWWYgVi1lLGO8x0r7jmPLDKzk2jOCItqs23VpoJ8
CCgSf0Dc6OSdAZUgCOPzRSvVabXudKWoz7KkqSctvJSFupbDFjUIgGF660/k8SR5n5KOfoQpWn4/
Mg6QU2lRfIi5+HDZAbUadvMe2zRqbZiK21qrB3DhKPHFR8tl3D2QrGbMF7hQO/xOKMFYJownHsCx
vY3AO1NFJoV587Ji5tcplRZ7HLrstEvjzvanPF5SuVq0YC28YMYWmrrTJOi0fJrNJTLldIIoTqbp
pj3u4VO576AI4n9IYw3deCy2DZOC6xIC5uehngVcVwRtNjLNcZ5qUNDzLQuNmTkg+3QPxatmfik0
AwCj4UdP/PZuTF8hvQpLGxqtIG9N6RcT6vnJHjAsokHTSMtav4Vt+UjESLqUALW8F6nhCwFSjwPT
EqUZBeo4qix2hr1QMh2ftXkmCjs8z/Mc60otEFbStn3wJW0vEV39/yntYN/H2Qh5hYYGHXl+3mrX
zd5dJQ3GZ9QKM2ro02LlNG99mmKlTwA89T2xqACK8NarMKOxCWiQc3YbfCjTeKx52s0WgRcLVZ2y
JVwU6hkdLNqP43ZBLfB6u8dV6ZEYvuwCD7lu5i5VFy6PEWY4Wrs+uaZ3iaP91Iwsup2H0JNJlYyX
YSHqNhaxjgXg/z4WOlj4Be9Sb9Q3CeZeOXZFH0rD+c6acalpOIBpS662LJNDCRs+VMt0kyuw7dAY
GFU6ZutEDkDHI99h5RK2xKiUuldD+YcOnYcRdwgrUAYumD0hN/dHkMd1sJJP/kBOlwlpJlwhT0Y8
4eSN1q7d8OLGZUmBl0NjDXWukI5j2ULe0ZQOebjzP9iojcLqIJRfQdoO1MW7xYys+Hg/UA0zIeHs
G7GSe6zFNlgPC6k4A9kgW8EsquDVi7zkxPQnFjuTnrX+omMw1gZrTrAW9gEJ8uizmsgVJlNtSbw2
yf2YBJ+6FuPgJW0IqAzmlL+t5Pqwvjz09S2dcZzwU/gj8CQXnhl6RKqMD1qXuQcP1+mY/s3/qZ5o
4vqIjfGMQIpgBS4YwsT9UlYEaS7a0MnI5Umq7tWnCTnhy1ue5Iwb5GhUsufGGquEwT+lL0p2yMPU
jlhR7ZSNcaX8swPeyXUAdgcMfw2VU4tJ4aa6lhBZioNuFZ1pfEf1nkKCebl42aNZ4bEMhZMMHMXd
12V+AmL2I6JncQ/HpBI91pdND6d+UM/89t85zMhK7+fUgQFPZmyazoDlDrFz8WxLvGYtbi2J8D01
uTpL8H8+mclQsGvCcd+54zIwr2NMrpVCveMqJ0OAsvvmzDcC6PjUesR6y7DS1ng1R0oFKRstGA1y
G2WRQLQIIN8Ok1ZKJcSGAe9Ek1/3NSbFderJRzc1kWmGBqhp1uiQH1rFqV36w2IvnoYrfccj7SBY
X0gyQtFMPQBkFWrORoYgQqO1t2mODHBipCr1W59LniWIw59Mvh8lgTNuvuo+ZKdykJLIj/IT37mj
KLawpdEcVCjtxGt4bxK6B45BTuSanBKe8iaz7hG4z5YxjS/ew28SXns+5M2hGW3Ljat43Aju52AS
bM2JEUWIti51PAUCePBi2GNewat6f9kpd42bGE8+aGmv6Hldc06NhD4nE2ogXbg8RAvsklBRDCQO
l5pQCHJPaz1Wx7C84htmIS0RSFI2g1dVw7iCMWsMAUPzi8yZUsoi4hRyihXYZyWZB4KQsQOA3E+5
0aa2C7L4UdGs6mZFPTJJJy6TtYiB2DsuQlaF+xETy7jM/ER+lfLPF6drfqbBnG0Ay5d6C+/TQgEu
OxitudtNlH0VUY1ZctKvn3OkYmu5JYanxMrsyZpuUpu9uI5Sh2OU5TM0GOCqb0gVmzvCfnLvjm7r
fb1Eaw2GZN94NKF1y3Pj2vp7mlg6eXMsOPKkISd5WIxV/HH9zi0DH6xlCL11SVqghX3LT9ZOU9Hx
XcLi517ALn0PjrMlrK3Vak4XqebuYL+p3orOwvcmNOt9+pYqXqW2AauZCpojf/DwAAoNQuNBU2Pn
RCVYOFHVeGuv5cjfXbu+FqThsSv/VuNokX/11Ut6G+XINiIMLKK945mxtFLd1BSvcze3PcjSHOl7
y0O+rQITbFo9XacG3ewuawK5dAZbzumizM8RXPEhDpG2IilNwzle0WNFH8dU7ZXCbJfaMmc6fApw
jS5nvA+Sn40Dr5t0Qiq+lK/sAhmwxPnMaPYMDffZaIWBcIdJtBhEDikwnpKT53or9oGS1dfnW837
vwE4uSVSkVz/D6C8nTG5tnaTm5JEQSUcM2rBRHyH3azW7TwsYjsKu3Gq2HfQfaafds7reJIuFDpL
cCdPPGOhhNM3izo5LvI+/vPNY829kR8UPSbRz6SK+9GAAeB3Rm0I0geezbqJUWsQ4VQ+z4L6JORC
A5qP6xLLMzd0JHEVYV4VrZxxBBXoEqta0nksW0fS21v3Nax0Db5NtPhDR88LLFPMEM0pnyCZYJ/d
cWO/Bq9M+DcmKGkZ3dmHvc2+WhwEv02sI0nPoVIMVG+kB+/9XtngY/enZNOhaXDhl4s66N5NHlHQ
F745efZA4maNxu8hEb2YHbuUW+CjUHb5YFNwicKLgoWzejJKqsvlFNgW+M4+yAGXYCLhBG4MpHe3
gzt/sEN865+5DNiHxMqkhfDz/Z52IUXz9bMuPzurC13JmGtfoiravekgOp/Ie7Pq1WJ9z/XFVnjD
5/lMH3uCMgLePXIIQXUbbz8aXSjI7xBxvJMmg5pFP7oA4xMvnyndJRKRz2/H3B98RvuTn+asoRDj
FWxmx2KeXtr2wJgO+11ssVTiy1BE9VDx9xsuiaHZEYXhAIHTBqTf8hBEpTjK2VMKSsNS6fKsbJCE
EI/Bd+HjZ5qLLc4PQPghSuAZMwGLZtwirtS1t3qbrdBOvomDJuYXEildMFj9YtQWzzugVAG3gwUl
oBz4msLGaPfhlkR+thSOS2oeP9/lIrDGf29Q095TZDDZpIi+wfRqm37NGzvHYxAzTEmNr4oBjQjc
INEUIAdmQjApX8Sm6ECFA1Zo9OOxOOOJlbWN09jNjRd19ctLc2UQcHSl/EfBVJXzQRn9O0EHVt1o
DfRx7uSwJdH8RrjoIMbgWDfS+tE/ATBaoA0lMY8Mn8lIZFy2yX5rjA1RA8HFM/EAfsDydUZT/HS3
1UHnE8oNqXJu4CGAidG0WQ0AV5KgAgai0cKxnf4Y7COKHcJLmPLSacT8dkF2h8Oq6hYBwl1oFEbO
bAnRO1X3L5+u3LRN4bZiNX4wOaW8r4BtJFJwj/G9u1fLTSuMaCx/ZA97Zsq/zU+jCA5M4jJiWpy0
skDSAXW3kgwXIoxkp9ScRpPDEnvchsYxOdZANqcJTGotCYsqJi7MWBL5C18/4bjsDG6zTEUvbr2Z
qFETsNXaj3LOnckVS+r6CKrGxvc5vWwXkdblk6oi5jAeFGsJ7Uo2iDRFKzowFDsqAA7xELfbEr0q
SeglnzMZ82jdvDfJvhTeMYA1t6g0Hcrujark9ORD/iHx6WopkK0rZiHGiYXfIUF1BZ4PBRVKaDSy
Y3MGZB0blll+WNoTk7VvK2/tIeWgu6qtergQBGBXUT1luxKGYoOviihtvhw098gDLoqSbZlYvQYk
T9pSuS1T0qQrBHE3PM4r8X46SkYWbSXYZiH1PvncZUVqy6mgRpW4l/9J+QCNKRU/nw6inu80f3Bm
eRlbsNkxSqnBFrvPeVoO5n/WaRrv1lYXxHj2wG/Xe8UmLqeyO7f/xRW8wlN1r0pK6vE3G39zxlQV
ENu3TKCV7qMt8QOJmUHL4PVIlgv9ucEzJJFgN0492pCsXjwFulN7Idp7qRbh9WmHr0UK4u5Q8HJ0
VBgkCAE/KipK3OEzzMwGeTJY6a14TWlFtNQgOHXySO4G0SMGU7lCrda/Tr0aByKJbVe7BnbVGKAy
hRQJpg0fWZ47xsFae5XErZUh31ZSjj7GMHuQY2qRZqxy7xBNZnqgqTlFeLFFd+ofCKFesrtBut99
x0vFFK+EIGe6qQedlgvZwxS45iDTn8fXIsHP9MjL4usUwH6Z5dCFtwiU23uQfHiJ2x5yUAyGLb+e
Z0jTQqXVCAqm2Wg1Rsf6xHyS5qRsocGbC6qFOPn1yRGYh5+aYMqVVPul45V33YM8kyX+IUEcR3p2
sfPKp3u3PP3h63T+RvcWpemBW+j1tfAdEEMUDMsFQAO3VD16VUvXwlj948vKsiIySdFWSsya7nwX
vMTx3/2WSnAG0o0BgmnAVFGBbExv60jX+D/R+ijasTgxnQ+ASN9D1nk/D7YLJEi3tU/DYNQyP/4P
rBOZGuix5t2B5LjnHjGsqD/2F1FZBudJ75E4cEBF4p5v/ZhQq3ai0gfHutP8WiQxmTf7DZRybcSv
1z7dwEyg+X+BZs2C/hUPBTLPeBjZN3xvVovb16xxAby055xlZ+UYwsfcPYw3GVM/YD5pb7Tp4//h
AXSkmCqqSW72MOpmTzVpWuoXz63kmp4S4apwWFvw2IWjl/pbr6VgT1+rYgFnblTDapN3BFZjbw0h
RoGyY809tHIqG9P5VL7kU+Wa8AlbUG/10mPApyCGx5TLkWrL7Ktj2ddTrmbtsV7rcGH/V6BiGUPb
RkAS5mxuvwYTutU291OF6c5ci4TQjnbAch767C9gN2n6Tb68mndxtmTGiGSD4+Ph3BSuDpCe67wr
DQA7Tg4WB88YKchU/6/XjFzZfH9akj6X66vVIDM5oxPSfrCivrzWbkQ8A0YXFpmLkWaeX+KU+gev
4xOnmD0MSDCgywE2dS8xL5nOIO2KzoaYsLG0fwLtFx6JnLTnhYUM/lVxz4qK4grqSJV6Na7tRkBT
vJNuk6IB+4H/JwZSzMLGL05YpdEcppW6DfGOIX9nqF+8TcbnYcPpHhXYhW0YyVRkdoVj9K4g9gRC
7L6mCTmPU2DmfyFPmoL5DvvCbJkdKNWeX0bfxh+/R0MbCURJH6+VPKkMGyXhtmo3UCUfLBVv/lgT
w9JeukuownicS2iwyaDx0YVEXApiRpy0E2jcidwmaAixMKu7OpA3BF6SXtoCZ80xLUCc0QHqfDLA
UPiciP6B+bltnYx2QoZpzlTym/GPC8eTduHab4tlTa1+iXw9gouLmdq/H4R8GOiEsPi7Mz02eruL
G6o27GZqnX5OwKDK9Am6MDcwFzYqqp/+up8Mrk+33BuzP8YdRHByH9tjTNCZPzecDcojsdlZBs7I
p6uYifLViSaDOp1uTO21op5kyo3kZS1AEOdu//+aORv0c5Ul38xuAYdzcizq05KYoTqCoWhPh/rQ
phQ8YLrHmyRToAmLY2BDTp0Z2I+RUts+wGBWwEgQQ6w92kSB8jaPe1VSbbCvFA6lDrzJ8jA/mDo6
tA1CB1XoOQhnv/fcoe719QYavGPHF+UOD6r5+cNRbSmWICigDch9fViSDB5/YvJASzInaQSU3xf1
t+LOFZEucztAIoMfesponqClafrUFN7BQf9zwTsIIQkMScLRDDG1USLRIhf2qkOrSTvfn1799HRC
mVo+wwt+0wTROWSLbiPune4aVe08dLbiq71o3lVya4q9bdsZW8aXY8qKcCILt38EZMMQ01uhNmlN
8LLfM2gt1Mhle5my9u5ew7rG84ZYV17YIebSfA7d2bzhKIHHoghereFEWbq5o/08xM4DrOhXmSnE
pzmoF3x34S0CDu8KBG4CcwdWTaAXYxwOAv58jkocV9dOy7+5APu+dUqQ2l1fC+d8LNX0Uao5tjnf
SbifT/IrLC8uUTieoo50ppHl5OihBkgWAVR7uhZnbem5/b0pAsj1YOc8b38RH0oh8hQhbpD7d4tg
eqQJmET5fiHmAjcJULR4mbx4frBX0xqn/46ff90Q7VJUuU/U8Ej4ofIM7wx3lfQZIX2E5M+mbPDS
CTnZeazz0EUeXa27Sq2SK+nQfob/btSPDesW+xM9wdZeX9lKeY5nXuh8aebegwAWxgi4n30yPqQ7
Puub159C+17p0bEMzBJB5UQ4Qj+q7P5aS+ddjT962XIKkZaehNX82AO2ur5iS+b1QsSoxWqAujOS
u8Qvp/DytKWdrEWdn69wnCk5CNMDT5evj8v6JI5oY8DGMjW4kY7RTN7zv5gwpuA1R6X8rjjBh3gi
ec4AiUSO+t0j46J6o2ui5UyMtgi8ezA64uZZksFEGYl3CNeu61kVyrQLl8Z1uuIfMR9zUxl9/ZYq
FiiuKy94CmUTce95Q6NaCxlmQIVn8KfNaPSJITAM4yr+PaCPJHyhS0OKsRfd1k1paHnXAOo5laqW
xfmZG50KtD3mVHnsLwPTuIHhl7oaK/Zg8tGQyc4CIfxrpa+Yi6npYCCmGbG8DtGfMrP4R4l3qpI2
tSlKA7bDH0FsuZJshcz7eYHK3sZT8moOeZT05qNHwLEcsFbhlHOWhRZ0I9VmInsGhQI1/O2uhi4z
7Z5CjvYTuSwsOd3ILQruZT7JIyw+ajsmU27AIbpwbj6DbdjD2eEaS9AnwWOLYm8P83u5hCJWefTK
z7YPoodUQ1gTrQxgE+gMrFOp6pg/jO4ymd4LoALjZY3fdFaw3WNHu57LH+M4IbV4EuFL9QK1Duxf
ZIU2xo7GlM06gbP5Yl/DdCxSQhuMTegZqIfY8Aeu+r8rk+HNRaYi3EwZLbm8YtvxMYOC7a8n01Kr
TLxcDABEGe7INfQY8kbnKguhj+pz/xzIHCuxULXHXHtQ3jshJnzqpuDMzqPRDnAqnbgtnmYxCsZG
nxclWFe0t7aj+GeJzEq6H+PAo80t8x2xVHKFFS597GLxbN8Y9QrX4ebiVvFELCih6OegxSn7QobZ
qAuCvb6Ze6FqBH5XvHXjG7G3J/Hq3e6hTa5x+PaCnnBNICh9PgE1hFvwVULoQ2CqsfQH3O5uMvu4
BJOLI8GrAgsI3bS2F7EQ3l9WeG1u6DKbRpluCUHD7Zn7OyNY23lEuDIGju33herR54Yu/Wq8+co/
2yzF4H+RJYDdkDmKfIcseGcsSO1xOHlGSBtRc6qt+iz9g/5t0SFcImgv/KWzQTmTmL7S5Gl/i2C8
/M9sso52pCMIVyCeliDrzK0z0GF+35xheYkozdle8UIiLUltR6j3NNz7K6CrZEb3BrupoThpMyZP
sdnpWQjrHUJ7WN1mfBomNWyn1taOrGGwXpud7nQoINkL0S/ND0l2uMgewoucKTyOqHo1I7jvikfs
m/USrCLm7PWOGTM4SCuGgLqLR4IlF6M2T+esnXkfIWS6PEFeDWSuL+1jjxxi7Re7DuNkB21SNaVA
pir4dRGKrazxgYqarpbjy2s/DyKzQjDT/nnOBECNImJ8VkBgP1YzqSaUAdljZGEjf28iVn3LEQGO
nzE5O36/dZDZadyZfzwVtrgf0ZwGen2u53Zv8vdhLj1oObcm2Fahr8DA6Pq93zD+4cHMkHM/dyzs
MgLe8MQV/iODuJcj8dwBEJQX65yrZhg9IVkOeWY84MYsA4KyLDpr8C1eZRBvm+eLh4q6MZfHpdnI
y+uqJ9avTpbS7buR924GmFm/8oxEcLb11v5S55ZDCgJkn6lS1uykr6sTT7+O7k0bptjgAf9s54vu
NsO4EFrYrlATepzu30Fc6+PXSPtGevZcfzbm7WazYgll00BCbLkv4Z/J3i5hb3ei3XanqGosK/yN
niPicNNgkPaCbiefyEXHT4WpITTtCjg0hKjzQ6plzthm8Wv/0ANqGZAfpGiWbPTL6Iti+NZftZbx
xWStVoufWAV7rlLn5tM7KsqkeOSso5Lybmr6XsGi1fu0CdCIio6AJ9JxKJ64YkVEzY+LED7gjYNA
GaHco47lSCkjoETxvnrsysk5irCy7mrI/DGxU9MyxhPz7DQT7FjLFzOlms6nCbLpnS3dUaoQVgZZ
ARyc3i0GRT4w7sDBxnYmxCWD5w6aUieJZjat474gwpbZgor8RcOFL/L9xVuDTNVA5Q+FcthERV9K
j9goc/OmJP55LpzBkX9yuq8vSRl9hg+nHnD6MHSOfx8tR4ipR3RQMfibxBv9/0gQ91bCEqPA0AW0
LOFRrZyZgW6ryQMmBXHoKyGQCRFOPepnWZhzTYd51p5ZqYwbA7QiV6S6kGJrNCzPo1/c/u2/ECDp
ZfSfVpKBb5PChBkkG0P1IhcIxIsvbjHRKkEM6TIFJOsHROdTGcJzSkPwVhginng6YnSFMcsKepYR
AO4Cyzg7xmc29Lo5ADeUFf7r6niO5a2qJmWzVSdE0IA76JLVh0ApHKD0ghVWFOdH9Dhkih30dMi6
3+qADRM0k9KObUv7NBVtPmWGIEPdvfCQ2hEDPnRolNSvGvLIYGslb507vw2fO6GoGXnOfzjI5Gxw
ied2PDCHR8wD40/TdBYS+DK3r0kNp+8pmlPgkQTcJxK1Oa8O6f+x4s/ti89BnHF2h/XIUquPGJgP
e4BOn3Twrvrs1E0PcSN+pc9FjSC1v4OkEegQLj89+sqVE/KAJ3dCrB7P3SSdtu8kTQWbldT7/3U7
HA1f+4pJ8sWIPX/h0YYNmYWPN6FR4o0ThlCdVyBcM8DHIpgx9AHYPjcrVA9QKNKECAHJlnM8x2U/
tMgIY/yIYMtHhRnOqn3Y1KcLYFdcPyerOe24Uiezcm75dscb69+wytN3DWxpU85sCsFl1hI83x29
kjUxKao2KKsAm///F1q2Ew4oaf01Jjmmf9i204kkiW7xdFs9b2hLDjJYQVm4easn3mAkR6wazsuB
6atj+gBBcGxcpEk9mkmT8H8eGwD/k4ActHqHCyY+DDTEy+/8XEfSw/FNCwo6uvYlicU1fwsiqeth
xOER4EEX+3O82SYj/xRfwcYOQQiW1ClIZlbwMtbD5+RNEJbbE5JqJwGv+9ojVh9ef+Kd0fAkJKF9
Db1NBNsynNkEYg1LGDUZq7Fe68/RC2+8WOXeL2L+FlnLjq9PSqInh02kzFVGmAqv0sr29BDaG8au
Mm+YnE6fnal8BxWygD01DfKzSI/oAgmgoWJrCQIqgFcO1wi2iq+AMi88PE8j5BWbkQvk4y9puhlw
x8kLO43qjV5u4c6PbKesPf9jnXgA2kDTz67PTjDpcp1rFFn+OKb781/XgR0V4NWwWLDuo/v/RFCi
n6lblSHBd6DRGzp5MIC1R9v2GXUEefNqz9LTxIdCW4UhigmfSBjhz/1cvz1H3TTAiLemmAc6NmXL
8LVSJPI5ExJTkI2DaMgirQ6/vSN5PziE58HG+AOiGQIHsO78lCSQYwPOGqxbeIbPc0Zm8IpKL8SQ
y7FE7WMSGjnK+bPcjx3QTmFKFcaEb9XtlxkulmN3bIyJyH/1WwbFB902/2oy0eBG5YwZMHonFRKb
WT2kIxDmlKLlRWGdgiDKz+EKOjBRnDx51lSg32ECLwclngCu+Xpl52c3gIDm7DLljDyjzt5N6dgj
ZJcLjJlg/mpNT0B52E7/ll5f/yROdbGKJdeKoCG4DGNqOcr7A4isCWGwkAfe/z/r8zIxHGdbx5OL
1Wd6iAAoPEk+/UkeFSgAIOGv/U8ThLluOztb6Rks4qwBmhqSK9BpW1GdGVQNf1wy86Xq10CNMKpQ
FVRwlO960evtE5tuMXWn4gj7FwVdhSJGDjOAXfDgxq9COvcarDT41ONUXANiXAjraKReVoZjKOYi
a0TPElCLxPNJX0In62gBQTLTAbPwt8ccwMtv1E9xK4xCu+zEzjm7d1e0CPeERkrY9eNVr4XjfCDh
TNm5+l+ErK2VolITheq4UAH4vCjRH0dhQ9VXZkCVrBm4X6F3bBMyVRq05k5K0XKeFmOvaKP2fwjD
rrdP5vZWOP9EGPvNpxuLI/RcamNB99lejjRpffuKvTBZsvvXdaCefCgUN4bZdHccjIwu62ehIkOM
xdriTxNjzBYGo+iiYdPJuGSYCrqoy/eSYLPrbgbQJYfnhgHEghR+UV2ICL0S6cEPu2WP0ttng5xk
ivuToEnDr4lr9C/uaIGb3iGD7BUY3NOYYHUYcDxUP3VT3KJFZopaqXTB+wqNfuueis0OL/CVUn8I
vOx2lFwQRFuPoPrbzLopMXgLtuwB6KIb/rqE0+wISKNJzyHEpsOTGqu7IibiaIF2ncFzbAHcjRW2
4rXy8EqOHuPWoaQvTgTz76HSI7fec6p5gI2agGzhDqfg86CnIcLnjz2XuzWbGUC/3k7TqfslEQEJ
2WdvNmSBhTPcbme8udz4O1CIBeFoDmYslgZDmbEFIRRY6zWGjZflvoUBIB+8VoCH1IDSjtda9w8O
IU8JjuLNBpWmiICENP9MZimvMa0w3B2DjLjTRpVXsdqCkJ7HWsZpJLJsi9Hk/VS318KvFKD2BxQb
F0uN8p1QoidC9qbtFPGB0T2CswOLQ+ZwBwr4FTilzV8t8EyJFLgFkBuRrfTE4Xjuk9FQ8Fjwpcef
lWpEQgAWOIGzUbPR6+/RtKw9NpLiJEd5JHj90Ezz0O9/dc7BYjqkEw4UtZ0JCV1u+2u2rQ1X//uy
iqZ3AcWRcHVUDq5gF7zUv9+CJqlMKPlBheYcLFX7Reo68dOqiS6/b3L5x6WOI/EBvEsT28pKtZAV
Ofg2DOyP9orkqCgmkRDJdsBEsmICsz+Z3+H1nfTm5KUWb+GqtUQTmrYMlGFAzTduzKsxuE5WBI/C
ficoUfk1welEFjtKZLhxcsEIc2zaMWWHVe6J8NiFSvodfF8RDLi5NKn94L2Yl9bjNrKGRBPWn09P
B6TlF1Fd9BK6PE/62keYBsodOWaUOXNMYinGPKt5Df+CkTSnWmfEVDh0mJSBD1B74aCAWrFYlG1v
WzeqxVMOBdmf9jOWmsNMOq2ndC9+p/yUB+y6NtwzSiB7P7BuYnxpv1BogImPkSg2czgdQWW4EQ8c
a8qqm+ddYo3GtWcC7bLBXaAYPQVxADzNzOJJBHtSVLbb1rxENWD1xEi3PC4jKES6e8b8xJBaKRPg
OWqRqbvk1bo22wYjsWm8+jwLF+FnZj2+85nIlyNrStHPo1QxuSyBSgyfPBMtlMckPKkqRXxmDJ09
mt/cFAPNNnhTgdgl247Xdy+2yLvnIf4qKXWfUSpcTehd/PD1YPOD83kzFiro1ti+WRyF3f4d9Lw9
NttLmR077ulJcE77aSgTOCbACoBzNYyI5mzPi7qQhRau+mu70ZCASoMdEknzmx9Cw03jSyVqt69E
/vbu+taQp0c+yuutkYoh4hiBW92ZN/TH8LstGZ38YpbZ6mQDGZJm5r7nUnKS9biy7SQ2n8TROEW3
J7r8Nude0eVIQSghjQRSox/f0PuIusu2e8eBLseD6a++1OhlJWBjkxAik75VGkBeNygGUtd27uJK
pwuP0GVKcE7YhNvX/eQaJZ4pd0Z7Ttxmsv4sMIe7CVIsel4SJNgwYe3Ud8z+y6EwfftpWHyR3S9d
Sg5tEHfj6etfxVcSCBU5HUxs9oZavGg8lXyKvkGP7zy+UAfDQH+lFtCdzAvVYW30OsND6SI44on/
1E9mHhZC5w0eYC1L66zwJzDSv8MWsqFvZqkeS/kP8SeZm2pf0BTO8jVP1lfSf9WeaKSKLIS0r9QC
u6VyCI3rDIUV3dB0BGNtEa7ttRDUPtx4SoZXCsV+LnwKICRgbzx9pfqjXN314+nCVp8hsdWf7SG/
zLJZ5ahSsHxk6XBmE9g3ws/fCpvg1Fg8qqW2u9coD8//YgkN4C34Ezmi8NltZROc7I/u7MZc6+di
vMJNZlC+vNF3Wj49/E11093KP+gXrsUzAPX9DiTQTXTCx/naQ1DST3uj0UD11Uy4uFtdig3WUflJ
wtizZ2oeI/g3uAR19fXIMRslbZHqBEc4DAisjBsyVd2Zmhc5/eFM0/2jJIcpcCGzWSoO1Qp884PA
R5w9TXtjTCzbxPlm3XIIMDNbr7fhj3H4wVUBGkeUJHcZmyUd7gfPgjptx3w2YwuQGDfbGuY1QNhl
TP21VVwcnsx39BHl2KaKkmpUIdUsbrEIJRGM16Fz/TIYUEgBCqwo+93p+lZLXbVfMK8yDoyLCvtZ
uY/FhYIfH4kAiPIgwF9ka54B/i54rJQxHmcxs11iuTVTugWwVuWmoauO8B8hRcc9teOPTGSbcn2c
IH1cJYZUI/WNeeqJqIWfIO2dcCRj9XRKAtO8Hu1dbkMebj5xBZkyx6y1dztEAKzDtTRhYhbCyQ1E
htvni5Tn1Q9qSNb+Ubg/JvUYox3G8SqUPmIS4YYtBBRQP7wu8F3JXqgl76/4A0/v2DBYe5puq4yO
O5IUDMWcTeVDay3ph3Z0AkDAMu6XNBXFBncdi9zkv3Agfpe4c76XHmcO+qfoEKeVH3OL2KXFbX2U
HCyDGqvrYnmuCkZUNndUl0FLmbC+p0somiOj2RxUoyHkk3yFHaMQTcbtXugg8VFHNU1JEAZvCH5Q
BVOY5MYqBn4Q8O9km5YHC8RS8Zme+/1BYKRAhy87em19elpxV34fqm6BBceOn624RYhFmdIZCmgh
g3CMz6lcBN3S6OqLvt1/ywEiT4+BcQ5TJWg1HJUGhs0HTI7zcj00JiaV2samOBi8l0tzEDLXx0Zz
gexg+xZJltw0N+SyQY/VlTB628YyCmBUKWF4dRtPjNehJuLkXjIiJ1Wm3LTBVPTBu3yrMWREasdj
peh2VE5pQlk9HnVWYaOprJfkI+60/6olt2MQJlpOYRym2PTsAG7ETIww6O9LvXMqAwJP3gMzyRpo
hxjAxc8DcMPiXkdsiEtL0M0CZLUyBYESnWiTuUo+Ub5IxIITn8UyZsDR6S5zf5ePUIjAg45DC46U
jAqA18LCmG6ewfnnovA2OYlzCEC1P48lbdTC3d04f9t4IpltOcdLBirZPKkKlVIgW1NnLdppClaW
HUIfWETFO6nXCWrQXMf9ylK9UYxXyQkXzZ4NAC5H1vFrdCwlKtuNWbLZJ7oNYv8lq0KA1sH0r+0X
46Ok+C201AwZnm3g8k8knApNbQHnLG+lbcq9jSIkDIOcip+qgko3jKzi5oKB+4mvEIgvQ/XPC+Bv
p1Kindx2WFNxEaNOmVrPamr74Xamm5vH/IpRHvGc9MN8/+GflH3pUtCUa4unkg+ZD5v5BGSPIxjL
hF1jjrrSi17QbySeN4TxqIcOTbeHM4t/9gsHtFKTCD4Lf9usEZW6WlcsV2BzKy40xuMLhrmT1tF0
XYM0k1q1ZiObJE2tKnbuTua4Nvpw2ItctmdXoqbBwVo+x6Fuz5td+Fn1N8cFOM5FqsdcHi7MehA4
GFiDzERIFf2K8CfEsEsh+2UFMX/O+UAP+K3Lz5Ov7Dezq7BwqvpRDZhw+qk7sQaQKKPNYItkTAol
NjEJJwQT/yaxxth/QCkWrmGRyxMX5Xs720HN96LlhmPTiirYR3PiClo0NlRfx1t9NGTMStZs8RPY
Vn1JOZzBZAYJ9w4Wx40K/28ccZMPT+HHf8C4mzqKEDPW5G9HMIYpXHufOj1YJSN/XmqcnB7ByoGY
RjOJYnUl+ZTKgSp0CYHkuADlRhfXKxCD7NlfJnahwVe2Qy0AdZ5V7LQXl733Ueo0q+bJJMRd1BVo
NkEEBqKboHzeO33KKFSXD/FurVQAmIntDdwKD8VONVOfiGtZYvCo3twLgzz5u9y6NGUcVZXAofmr
Xb3t8kEta/SjrSgNc4gc0nGkivZtG63XjvL1D5XL+FiO8J/DY/izPx7xMPe/aTVASY58pCEIJBPn
2dC29hhOzEMeI8iRWOFB3SHPLOwpH7VTwbtoka0n3JJptMAynMtJTyaycLTeEmHxSTjyzto/Bvi+
SpggxECOKfTA1KYn9Lfma+QpAH8fgkOEH+U9oETConkjO17C889Q+uBEJDQm5y/8JSWRucArISOR
/r+Rig2GmCamlK9LoPPohamQ7v9h3ztigeXUUKp4w8EgLwJ3DKgZglH+fBCdV3LLaKPnu1oBCZ1L
fiPkbjYKR0UlYjuXkRPWpbmUQYlA9vSlxlEPQaXfwUVoMhpj2WNxR2TeOtRa9mwwC9pgFWoZc7ck
uk6I0YBBwxzeR7M58vV43dqw+qDm3K1Zt/43dXBcj17058LkEOWdJqWaFemA2Qq44wh5mCHpGxo4
7NUa8CDYBYJuQR9b8dUPNt1FsIkdMRZMy5W4kcXLtL5njrJvlHClsGmHwPjuCe6BhVD/Q2EzbQdp
vHMk5x/vgNVzQ2snLS2VbBKat3VFwjkJ9intNULqcPVF2famDDhf3cQLjz3VYVqRW2xbpp8wbby4
WEYYiO+Eie0K/VTGMzXX9jpplEaLBIKgot33nqTqMOE5ziatCdps9iGi8EwT/UITHwbf2GfCgTe6
DH8vkqvkf5Nqq9AHsWXE49zQLqfETMrtMNYVMDqCokldcX7Mv6q6GE5CTDXo6B5p7SLACOyYIWgy
0cHiCWFEizDQRzS6oX12v79ehSC9Cct2YepE+za43DkY7SrIlhMzDg5JglUAG0Ft6VcGe9W6hKTD
pBF6ufySjyTguBAhuqZZonlTUDqjUN1qrtcyGVn1tZvk1W6Q91QWgPRwbdZUpIscOlUeePP5Vl/7
lsqnss2uxW7WIXSnGmBAeErs654/Et+QqwdQaiNOeB6PPy5pJHV+woSTQR+HexcR5HCF8XSo4ks2
DpPqx5iGAi4cYUJOmzn9FYRuzndGfr4vnEqeAok4aAIiKO9GbMmnD5lTd2oC7/MloRc42izlj0WA
KCeiory6qwcyK4p1qSXz6S8Ixzhdh1UAY1mEZFV5IUsDyugA1hDI4xgEFeGKP0De06/oNN0wJcye
yON5MZlDWRURCs8SWEhlEcFdAJ7L0Qo6DvC8VvL8MSY8nEoXEOweo1Y2liBmMV42hpCoUuP1PwZk
mt6rRCe/tsvc3jOcShPklWXtcvH0TTv0fEg+Z8h2PSoubZplP6yFvs5SbDGax424nFshI/pkUEP5
cjulBs6QSfQ8+y9wls0/JvoXQNzmmRlvUfARAzafCMSVwdo6bfFS3olpUvFCMTnHquxs4flv+1It
5ved236LwOCs71EdhxYd5mltzRLIvlYLLJDGyt7fxLwRy8ddFnYhiJ8wA9gwAHQFBhZR/G3a5moV
I2A1F1SNjlADUZoZ4/ow0AShfW95ERi5W3uSIRVGy2Kbn9u5k+W9o7mDL7FvDgsa/wxy5m8v+tiK
0+RGsgPYN9JMM85S66htWT8yLqmHJ2CeUYL7VScvpISNA8IdJ3IjQUrWr2XcNMHWZe7GmxQicf8B
TkV6AZmUZZ7Yt5Oarx9xIu1KhkOfBAKgnvx+5Da0us306sQqQHt0Lu4hGMTkFZOzKEllWlBm+kTg
qxCbUneSWLUArHtk+ZRBhI2OlVcMBjg0P5ZrxbxSgbkOo9bJyzXvsNQ4YOVHnEP7FxHQlQfsGA8l
GCJzn/Rpk4V2WBOFdePqw2BJp9iobm5vPTt8TLROgdOYq5z1787qunFbjwAQH9RVTzL4RHqJSW/j
Fzr2OjQPwnCW4Nmh2zWlaskg2vAkFa4WAr+VChWLV4qYJ0Ewx5hS9SZdv/mqrA63ecxxiZnozLd4
wCiIzoVvyi/0qCiHdvFFTd9fzsDvfqkb+4DZJdMMrRgosXDhf4IC990mLvJwe+M+zioGlI4ybG5D
oOlVb2TxdNYKA9Fx1SmImvM8Gm+YtilDwJg9qqpazTztCSxfF4jB7BeSAtoUCh8RXIPNC/ayl1tP
NW9kYCnsW06FIVuoTdBMqiOkuq2K+PpfN3youWmyFAo+Uo6dIdhfOvXlouDFxcsV2tli3Tvjccft
6JpMo4QxzkSojhCxwYS1RnJXtchYPD+4jDvhQ7iJ/ogL0xo//HEBEe9JGj/VCXWr+o1NyfM1m6Da
ltfGUtHwMkdLtGqd+JNqjGTSeEdcXX3DL5LU9dXVUBWxTdnRLLltDG3jsBjqlo/SC3MjOWjGdxEc
pivTbzv6iTZoz93uGMhUllDqHxp1o7ooHL2h4pxE7yE2BAQ2Z4duIxBVpx2o0pjH5zeb2iywdzob
YDhm4HKIQRsvWDAaLIkLGcv67HvVLGf9vzvy9BDXjVenXshsWPt7HEi6QxqWb7fz96kwAHIlW8sy
k12dlksBjSN+4RabJikHQ4gyI3tLdkeyGzysSxJk10dj0XX5gVUAL0DJPXymz6HZHJRzUCZiRgyX
oERZLTKuzqflLl2NgiWQEDIOx3Fr8uNTu48tIyC9IQc+gtOQNVtqopu168FyE4iH3X0Mx9I0sjA7
wuEC6VBzr1EytU2DULWTVo5b8IunnPq2nbp1Ki0WB/LaR2DqXNUvWhLRRLLUQouqTa+SgmW2EHXo
pD2MHlOjKsRSvPMRHpHp/V/wKeSv9Xi7pc/obVpsbJU1/d0XTyxDjh0CNveAUzPx1r62kA6teJI4
vd9soLZcnKIyN9sxfVsNYV51nUjNOEi3je++qnoz8nW+l1Xs7VjQ8eXy37APbobzAITMFJISOOD8
7MA7gK0YjQF4TNXZsf95XEYjubL/t93OEc3mtEyTT0oxS4zFZJcHWJh0+0Rca/EcTb4eBH9YeGSa
XCidjpO01X841F30Zogm68dXbDQ5TzS4qxllr711VEyxoPVW4xtV1xOquxOWYoVl/JARBw/xPTRd
P74BfDEe/Wn2CvAIbP/Kyd2GCJ7Cm0Ep/CqmwdfyWaZ8IjZldfuhteVG8KSfQuzEl2fjIe6Etmh8
yIKakTkcrubgfEJURTpBpA6DB/OWalWhPwJdaX6ZyuVZDaDeH9fzSjZp7m0kvXmVPrYIIZ0gFxUP
CzoGGuEIDgEjHdjkHijyPSIw+fCcKwFAGP2SSF3funOGf7scXeWJen9lg9JIFVJc7ZwJzdlzEZkt
PYDr/tHOGrpWlRjROn/L2IEpMwGKkVJJ5sLjDQrkF0IC/2xPd+j4FFsAPeLTdGQfsUSs4hXT4+vI
zA/txdZkxZtkVjErvAvNtOBptuds5ieQDoxnSgAvyfZcQMdDyqDS9AoXsyenOUM1Ik9IzTJ1iaqQ
GkewEXqiOQ2jxNnkKLhEBvLrK9hsSm/fbhbSEnj56DeaNZnx08NnKdmH8tDGrS+S0urXDQewkPXf
ZU7WoBLX/nAqo6jzpFMPxNxSvUjjDFQLr2G4T2KjSsjlnn57lw82XrVmJn4Qp5GiDZDjDt0DiKNe
Pe55x9oxVwwo0hHZlTO4Bo7mcb2NpWL/FmnJ54WM1l7H148fmKHE4QuX+D7WBPklDk0nJ4ptw0gG
CcmfCxgrNzmYG7ZuJnqUP1sw1gv5f5cjwE2H5CWWIk3/jM/OQMvGppwGq2xqftqjuiD8dJf2A+MU
SJPDylnPYw8N6Nvsvm4elRKFN80TMTIb7z5i4jrWu7QSNl/xsMql7LuKnYXJ0IWf48h9cpgXF8JM
9NtI+NnoB6wfxFAOCJvp+7ZXRjs3nqHP7ZNKUL4iofAIrSDkYKn09YOS0aWZ4DG7QsyjfxB6ANK0
6dfABhs2kI39wjt7Yo1Z0K3toqw45xFEsAGc23hHgcJG0vD0sMtjzv7TMeXWPzJJ+/ew2AmP84Kp
s+QIY+o6vDNPcUs1BWZoakTWGeWNcgE3m7T3z+k4s/KSojyGjh2z6rvqopbuVolDtmvB6kXoluch
xXlG2ihQCCunAaAjPc1HjiX1Ef27Qm4aHhYVYKuW2Y+OtKT5sB8P0YKuLpTrnVccgLzvB/B4DR5X
NEgM8ygOh3G53LpnRKss4IGadL+ZGTBAiMQYZNtsybY1x6nWTIQNKMcAdJ4eJGqzvdasHqMrTPQi
T61QuPWu0YvipkdlxC67NpexDhrZJ3G0ERYyQ4ZS8QzifeLf8f9Qjrefm+9XuSwZaJIFElAXogut
8oLtcxZ5/2gl64UPoNruEA2/5xc1FoSsZlN8ylYcxgzbEc2KMw7okXds93K1pr6fajU7zeUkpDdM
rsfHhAt7Sxr4swjH6EGN9ONG5PMx1aTBKT3+GmtRqwGHFfwCcXGbuyo5wQ88irRAG0To9bA6m3Yj
Kjl2hsEiEqdOxW7cwG2xTW1Pw/cJ2T098P3CHT2Z1avByPud3e6A7H3RxVYdY5XcHvcK/gUd7e3q
RPg+k879WCrMLm0G3MUscLcootX0GeGscGjam2kgg/ve1NEmvF7zVn1zkyN5McT6nF+zTLkls5Rs
LIlRxpztXUoqrHdbOyvdsIT6mYnxZ+Qad04/wDNWxIKhOY8N2VuaBAlG5OWN/VmGXgi1xNdb45wd
ycSOohDsbl6FzjN/h8U/oRCY29bGiXMh6FyP8DUyfsPlRN/KXTUhWt8eA08Bzzq3nsvw8CYi6Zqp
xBsSt4MksBt7AjgvWb7QG5LZ5Ksbvsyc3jrTXXBAAqf8U6MwUvdArKb2zph7O/cAfOInuJdXp9WI
gL1NUr2F6iCKEriyzgEmEruZcryd+qY+z6A+Vm2i3HFWsOgHC9fuaJsZlvRnAkAmu90AzIpvnSZ2
oZWZkqmIlGhmiH6WN66dWcSLTu0ucX/Qhh2Atqym9tUn+27wlWVRG1n2YH5tRiM8y2LnIukv3MEd
ILQkg796fxbOZsTfYQaNssk3UjTV6vLfxv2Logp485pInPZ6UwLFMkvNnB751Y5hDZG3SXCswXv0
myZpkLkK6g7wdyCLs5aQXFZYbdy/no4hkD85/ISLH2pbnmCRW5nDtWKmvI5EGDHc3LL3pUoPYwZp
at3bNo22puN6yCYQ52dtUxdvTBqAngTqrpdUDU3rt+X99vw+ecgbWvK4aK/YLhotGBHKl5fMOF8e
5qkXKh93pLhf60xg4LUd9pIG147I4vGqk4eRE9/pkqgeuA/g6QW1+MUeme/9Mcocp5CpwQ5lBg31
WTfbBrO9ked/RcnL9PLInXIT2A2gjZIpKEXZp4EsHRefvuhuvJlWZawIAkNWK83tb/li2IhJPdP0
1T/vc/fkCNWObGczdkCIAMRgseyrfeB4pGe+EFdYcKf1iXLc79U5y3hHEnDyBBtAnT6xFsM5rQcg
T+S4V+HlU3O3SgUbJAWktu1UWoh3G9qDH+dXcBdCD0Bxhj90NbAiS+ZqphOPUKQWZpvckzKOeO8n
TjqhufuJTnb4LH/UTPtUzXO6BOrepedXXq+4lcg0ZYUQ/E+nGA7enk9pUwefTsrn8dpCilUfB4GF
rbk5FDqgHIMpnV6LPwnjWmncMNuouSPUqP8owEGheM2XOLPBTs/WuYND/+BatVvEi/1IJXsJNlN0
+ebju/49YM5QVy/EKEshpW9CjnzmGWiu/u7cf0jCIA9pzqVC0pV+P6jcP0lQb6JPIS22kOOTadEB
RZ/OcZ8JXps9OcyKnNRdZUscePbbjAOQE6NMfvC16GWB8rfzaoZ7VKibi2A862oFBHrBykqSTRbH
gglVeF+CrvvUoovDLizh/MOwpRkW2f5Ruk/3soZtmQX32BnlaWH46qcyqtuhiwjAd0YuxlCivBlS
Mn1TRW1bCkaNMbZYFz5j3ZJdXGafSswgqyctfI9Tx9EaEW6adjtzPeFWPzGX1HCFjAicyTM/A41J
x9tThjPAp+/1JX6fWaNU4HsDYxPfTrbPn5F1r/m4uA/lJNfup/sRt5g4Dwm2ND2hT5UTrX4k5bQY
AXeX96ubQR+y1fSqEE7I9ZYOm91bptPeV1qVBmOFSiTgw7FJx4qhv1CPnyvU6dxI3lEKwe6N1Z4j
t003OlG/BVhGhaGqRMpdKbrCF58DAEAUJ8h7Q1WmIcK6NCchgbxjS2nzrbPj0QBw/UwB5TM0U/4b
FqDsXAbNbritGpSW+usf73bTP4wyyTbGLOWdRGcMLtdHzAgLOoYg8RgSQPQEwQHSewhSp0sbM9XB
6HzMMoGhviSATtmC58t9dzz672z3JyEgUfw1zLSGxRBkE7jhQWFPU7LQ5yqTjMmZL/pgQkM/TX4V
Viy3pLMhc037wVOO7uQTe6oictUJx7hOQ9Op8LMkSLQvs4r9xBcn+CaQXk9GVPmxU6sc9YFW6cOF
mVrOGlqzVyRCKUQgn6dqU5v8ht9V/pE6JJvE/q9ELn4dCwIIV1UObVxkhIryY8YE9WnSmCHbnJuX
8pl7CKEd9G8HLuXFDy7a6NZzRdOxpYyLTN+womOUXkkvI55ZmFse7kDQjUBcdcgIAGOCgvU694+X
rpa/ZY1I7mM8B50dfktdGiJ5//i3hlfovuZvM9NZXWy1tvg913aSEN2AAQAaARRM5IWw4e7i8Chn
pvG/TNeTb0uemdo0bL7dsAzVQ4L9ii5RDyCmrKAdt6F+KIL7AMhrYcm/5bMkX4iw4PhDEwIFoDJm
UqsMeQBmznLsGw7xnmwsfiNFXS5NQy/TdqI44+zjU5bo6Vr6LFoJyPzGm9mIOCpr17lUd0RdzrlC
1I8ykmm961S18CjWPondC8LRulm3oTJcsRxvePbvToB2r/UVC2bByTVvKc8yHO9GspLUvtU6H3bO
YzJZ3v20Kpu3r4i/IhHa/lIEdRrmBwKWRg8U7MjI2fLOzK3eTRFiVsStfTVAHolomVhP1KXt/fs7
PF6SXSmE8nyhgvmPkAM2zAwvaDOXY0zX50YK8YLLzJ3mTe2zLUmk/PE+neuMLWjeZf+ubggnYUoN
CjBDstCrLbEQ88FWh6sGnOSeyR8qVrfzuJ5CTlB7U5R+haJnZU/mIDySZIu/ZChiEsTuRnTGhEN8
VjsGpXT7Wy2R6vJ96aXnYjCMVOxWTozigdvGYwv+G/9+P3WRAuiVRsJES5jtOAA4PiHFM2wCZSIk
x1Uxz3B72id/4q1CXsrjk7ddhvZUd7/4yTUtBuYLr5S+obxKSdW08l6u0IKTkw+ZC1iM8IeciacX
cHmvcTYUgqCmNrRtF/oYmnrKhA2cG46c0pKZdkxPBmXLcJnQLx8jGt5k9ZSXctxNj5iISOgsiypQ
qmCFCD4Q8Ax/wlpBKXjGs8rX58YaKzOHgGukbIiJ2fbVqbPacJTAmv0GkHjpiHQClUs6zFzIAh0p
xfZsKzOz40Go14VrGgVgZiRNdL1BUU+AA1Ci0P46oeaMNUIyWYlC5RXdXnOjzJIiz2tpPjLymzOw
Es10OkX1I35ouKmH6rs69sODIyLJEHSXzmdTLI/8P2O7boqmGQCwmHg+tU6PyZhPFRsfaRDDJpjt
wsomEBXFb4TrdSqpTV9eUVrfEMbt0o5zImbRhl8us7rNW+sxhYNvmVFbI56gnPXMaN/FY3sbzKco
uJ/xrgu2v/jiJChw36kd5DE18xtvLo7Vlxkeh35QEI235S92SxIujUhqCUApy+eP7SFZkKhtjyaK
4lFEnaHK9V2MwoA31dfVGrxp/Gli0B6ZD5NAQ2iJNMKqhJFiXg3RW/ZpyKDqX1R0pt71fJoYFFQS
09Rtz0/9gcPw01ZjVJxpYPKF20bRIQoSzPStKj6M2nVYsHQ58G0vVJPru208KccKUTHMqjmHr2uj
Ykz5m661apHGyrPGuXQydnKPqMT3uGkRDPUPxfNrQeBVBMmP4hO+6Yv6JbrPdQYskV3n0bddb7Ui
em5IQlNRfj+LeX/wYdjvKQ9LXwnqoda84VC5seCw52JO0uLWLMnk4mu4VasNZwiVXvpvohpnm9db
SYeKoDa8MLtJtd3Vk8FdAkk+OMyONuvxSWPkVkjYP6pCcK4LP83cY8jM9X/WzLNRmNcMs+L6i0e4
lZm4P9T9dI1ePd++4UFhm/BQfhIHnpvrHppRd5BM9l1Qw7hp95ma4ZyY+BK0tzL4nNvo1Fou8yrF
JLDDaKQVmSou8UxdUjrQ5roDhgGIqYUGyXdTBNJxYMbYD+6Ju1XbmnoYWaimt5FZQLSgnyzoy39t
Kudk8uoPHCjtlKqejeCqV+Vt/i3YChbMuXeZy+IBzG+ye93EuWyEPU+WaLJq3lQyn9ZehaCDPHBY
bJS+JqJDf/b+MoQhF82eGC0enkJ+eMjpzuk4GEQ9UGuruzIj+w6cfDya0l0TA2aumVrFPymVrOOo
TEeuJ770d7a1MuAKh3D70jXF3IF5yJvznEKtMQQCBAbyKamom6p+ALCa00LHWDDepk1o9Py5Dz3Y
7gLhaW1ydoxD/btndj83ZGfAbR+rJARo0QvWMUmssIYPpmUVgIFWjlw1gbn/yt6iu+5A9ChaKzRo
q0DfYY4vEVA0ZQshU7ng3UhyD37nQ/9GIerPsVeqnDevoyMGpEJdx+iuHq9A2n/8Cae4RKymfvMp
7bjPaO/Zeoi5uu9MtrMhxYwrLHBdyZ/6Ccpr9b1/dZIMY2GLGGkn0XLhTCyUGbNUrGhBR6Bdp/Fn
UgAq1RVRQJ4j7eUzysNw5SrwD9EiiV+5xQDEsPQAIAh9w54Bix4UWwRWc+DA4L5r52x/tz4dQ4WK
EpP4zc2GeZ3W7Q6spGWjyfTGBUVYlbhnZSF1asQIA7k1fZV5y5Eo/8lcZbNJr0nPuMWq9vdIkLcI
F5f2A3HmeBJ3rprCsP6/wqShoCKqftEbFafovBpMMMRpI2/raiwps5IKK4CNqFLcL0gS93nLg/Ys
ONdO7HBA6tORLQuJ8LlWWXb3CXZ8fFUMlA1AV9nIgBJKH+pUBkGjQtyJ6q4zkl7NVsS6vUKHEdVE
312P7wtdU9KigqkuzdI/poWiznNLnKEiLU8T71bfrh4KEer7++Ougt6AfZSof5ErVAFECTcaqQOR
W40PAJyO7rZNYS72EYian4FE5GnfDnmUFrd+c0Wj3gb9+42rsrbu4UvhU8UTduSC/bGIopr2zxOW
Tj3dROkLDsklfDkFdkbx7m2ga9cAIFvYo/NgWl3TuffhFzwOLjUYirNqiug5EkZ5URsFsA6fKQXt
xuzIN94NahaEvpBEULzRft9dShN67NBBgkkeNisd62XsyxEHCeRSqzTaVePPZmA9l0lRhRTAy/L+
CgTlVWath06P0ABhN9C/J9vZq0Z4/H8pnHn1zSL9Cuz64QVFA2eVNNCEiXlxi9dvCAeCzqZfeSLL
ePVBTEBbYKyPZzW5a/TEcKeFzc5wvjMj7wj3Kcxzwxw6bfe6+FasY54nmSqqufAk7Hwvh2JCjMNZ
ci6GrLaMj53oxSyULpWzQwprfAmoN9gozf97rQKbBqYjWKWyQ/x78/tW1xGzQ5vYcRwWyph7Mr0e
xkbzmPX8z4hS1HU5SSA9WSVvUkcrUP3zYmtnNhCIw1/LfwhofS75EPEAGAaCsaEMfd+cQQ+esTRn
PeLyYII6wHwGbVqd7sZuL2xSI4udWob/v6Zv6yJXA45wOikVmWgiZpWzZtKuGQw618aILEpHXyeK
92gHrjmkuO2MRECiwTlOpDxzDNCOETSCoLUcPFW+I3FyfmYtOyu3PuACoIox7rn6hNeELk0efzkl
hQJCAJDcTyUdqm6KExMYXxjChK0NTYyAxkittfQyRsLRkybElCfV+OuKVfosUIJwKtLC1+sj2Mv/
+YmmmiHLJuyNGFA//e39GKcWiriqjWbY9YxByihSHqrZxYmCUnRC1cNea8y5tmILp2vdo1D1YN9q
ay4tXJzybKIq8f0067c6p0Q9aAb1YyVN3HHhNWWV/gjoO32yvo5XsQ6Di2QfZ1WH7ixcRabjJmeb
3vqX1r+h/Usw60+ad/US2dVER1CQho0Vt87M1KLjEQin9Fyc1rtAOxSGcbzdhSY0lCnVrxPFzILY
ESPcbeYjN30fdMTvWaoLT9Z06Z7EpNyrG2aokmKuntAI73UT4J0DQx5sopiT9UpGzqtdyzyFzcZ2
I8y9k3lGq2xPSed8TFYhy6qEGRaLbgVZCJSzZEY0AxHxVe9n8gBLZsOwW0AFpjYJy4j9gBea1DWZ
KHj68Cx8eEeL+hoJSMdRdoz8EwBEz6tpKB1fMb9P/fzbfwQFXooCfI37Jbi9aVACrsDBCcFzMHw0
vcqnXnLJGI6Kb9iA6/MjZAe3INYF4k3yeFhyWqMvHu1IsY8e+a4rXNo3wI1ewB7PgFJhuubxAYor
mVhidknhRsILvF5akJ1+xUxlf3/GdZKX0SE+jkGtoqEnDMnvLemmZ1oejZjI7yclFQ0Tv3UOk9g5
Apmu/afE2kqxZulXBA+1wwhfk7bBW+Dw4H55bufACQ1zPL1ncZ5NVBC1Fltodez2GGGmc5aDfeGS
uUlge4f8HsAe8QFs9HQf6e7F5hWxgSEGJVRLlbXvAn1rR/Uje0Wsat0hqPBdgNS1tWI0hFCT5HVt
xquKF+CiPvREX76H+xHlwMhGQ0W3Kk2d55eEgu2t2KRIKtG41KVrYT87Eiqi6w07TPUSmMtudqnP
MMk48mDB5/r5SvLl7mZ4uldbdAmZTuDMJVdgQtshJCsjD91WzdHcAj203rAoJpQHkQdCEctCxtix
S8Sv1q4Vze+QFUVmI1gj38xUiVDSRM1PG6FsZXds87Mjb0+FNXwhbT29wQuhdTge6qP9eHZt9IUn
gzRCvh/Mn1s3BKCgp6vYEVGu773WkRrgs/LnFgNaIc1Zmo4LWYK1PXKrTA6G9HiJfDNVZaxL7F7s
i54DXA28iSUUQZkBk2i8jjPWNxDRInwh7ZbnWFREKgThWDopUZMRIyeaMRC2/R299TxeU5FBrOCk
kf/Q27J8lrLSOygAVIrMNHSLVZ8LqDhjf38A6TJPXLh//FANBZG3OG/ylhENKeBtrhDqV5EybFXZ
beAK1Df0+LNFNpD5hdh42k66Fl9wO7WUpL+kpyUOk7HnxNva41hJQtw9OdN3xKYCaFvxjJ1IRNSe
TnFzUXg/4UKc03UAZm/UKc8qf9xiStyqjWOU9LX2EaAF+3XcbURaWgK0QCtrdTfE8E+ccGdFI+6j
eVHfJWeF+/VgzUQ5Hv/nTNbAaDH0cVupXas53taewR0HfZpS37BHSagH0MnVy3JSqTYCRI2gJKvb
Jw3ycBnjbG0vtyBNWbQWBd/xZkpCN9AxEMjghRiefltQuXEXUsKcnTsz+5BkOpfwR8HdceUzUagF
Gl7qkZocf0YUqk01bhmhIjWUQVxhltmUBxHEbY6t043UaXGQk/5He9O0oRp1Fd4Ktcwwwg9DMGpd
wTq7rxFacxlIFVTw3ZrQDJB9Lt4rzRmyMt0VoNIw/VNNrDglMvh3gwR6dm1gDSrfVZu2/VXQhjtI
kucIjl0UNOZMKNoVO77ao1JXSjvtHo8F4/LcrBaeDdB6b3O4S9pFki07JKIynnZfupf9o4renm7Q
8Eqjyna27UE2b33MNP3sso00rwRnRmJaAbRrdV5Z1BJNPSq5SWA8mNsuKlcHqNAzNEN13IXmdV9X
ofJqNqBcciXGR4sKROieHOsfhcHJHAQ2YN37/pxIM2XHyNOc+L+DmJ3GQRML546Nld18sJPg9D48
8Ze8eJa8iszlTJfCgl7PSuN2BIAtRl3WOcDnz4ZW2pnn5ZJR/LKJcnhPLzSC5BWbnPc6zClZFw5b
kxIjeNvsIVuXI8/WH2B7sIUZHHzcfgsbckPhq7qRkudzSDSkgq3XrWqLZGAon7vHk4HDPXf02z/k
3N3siVj6adNQ5t7dkZpp9t79fzBbO+TC8/tZPA+wY+D9S4/nqfhhPSSCfbQbEcKQTFOeyXoJHgYb
FAoYRcIUKCPenwsdN819HyV+37TxZ0SfB3+Gb39WrtIamb5c+dvwQS0LyY8ND0nQ2uNv2EVZpXVW
vXFTDmfFAe5n3Gb9C6e/7F1WdC0qPzJyA9zN7YXJ9ZSg8mMW6ECtAjK/phbo7wTAYuONO1xslPTs
nMimeAEWtYEvWY0FsM2ABTv8eW3Gp9NQzMi4Ydc7lQaKaOwNvjyq3IilLSV+uUbgHqrnP4apc7r1
D5+jMVZ2nz1gUc89knE8cABzW5CzT3uetG01tOy9ocins0ZA2DNnqZmonJWAg3AWGVtcmUs+zq4D
/j4RWZePBk0KC07QFCt8x/s15AHIOvIfFPAJpeNg/FUyKos9RWXh3wcuSW9SlGeXgXYQoFmR5v88
/TSQSkokwBhFkvWNvZuqF1KV6JzzhscJSDq390ZmtiBItXOOQUCtZBoQy+1mQSfvCkF0BpHMbGGQ
4VyFaAaYDgeQrbSx7e9pIBl0iomjEEig3yEhn3G8ftfW9bsD0ygl5+15Sgi5rRWd8mB83HICmp7Y
ldEYpcXy2iw4dgHGWIfu7/0cpqSfiGSIGJn3ElLIowU3uzD1k5sLyz6mk175wN8+Ng6HfeUSnKRu
r63EHcQ97ryA3m0OdWmizxDJCkoVNwiWTj7Xgv0KgCVfB4XUyzOUQujSEue9Q61p2UVfaQsqaJQQ
5u2Yt7Tfabq7eV0CYYGG+us7F0ccvY7Kg3MgPiWCGE5iGNJLXqjmriKJsxcIKhQhufrrz0ODx8v9
YD4rYQMSYbxwlDokJtRtyUfLhOTnmEeR1dHSgezXrcF93vL02FIbRQouz7A3pXs0v2/QsW4PY+oX
nXLWpmihWrXaeldMJ4A4Bb/wgxcrN6/cgH+igjmzHPnK2rN2TG+ZDDQgrGgiConnITsbchoeDt1i
RHFp8VAK1VSZFvmgW6dzEq11JdEAT9tIiDte0XFv0EQ1bwHhJC3c5XoKjweTH1vuwlt8BLBPzrSC
NNDgV3jfm2tS1WQvAToYUelazk1CNJMU+ZL3f3d0NkMcJP8OjITgTkEX34WmXM/qgjBQIxHYsGZf
TJuQhQ9x+GAfbg38beQOoWaXCtatZn1kT8xjYtYtfZMwBeMEZWsB6i37QnSsiDH4f8FGLebEaM5t
v8hEzo6kxxcvAnGn1OTVaryK8uU4fHY7burrfoEu0NxVibFgQCP8H+0vihM5nBtZtvqChTdwff7r
sq7Qm+KTl9BsxcEolGp/SWktL5rzzSgjVmbQtgAuRKwDPrv76QS5V8/HmW9PCIc7LhN5vgPIwDJq
BRSVFPI1XKH4NohuEimmfGmRDVohElrOV8LNmRRawvnr51ziglECcQokKcAR8forW+mJIMVWQY8A
+m2N88xhgtb/tcop2Lm/6Uv54KwDj9kfIZ8PdXOB21FpERfY4GoEFJMuc6ajBRjBmP1AFMGBA12D
GzjhaPadVqzOLAZpsNXnJLgHlVGo9NSupKJmoJPg7AIJSzAImUjhsc/fnr7JEKSuqiVxH/VqNUQl
gdPQjDngXpKP8sFuWpUSO4eE0uqPPr2MeWW9X3lExGfWzntXtL3s/rRYK5LTbK3OlfkE2xZwHpgZ
HGQ65kxcaRaw6RndQRl9xkthwhhS+kAl+AMntoY4xrqraum28mLPGAmAVb9lTJq2nUBRb7b7E7hg
iGYB4BdDsUZVN7675YvsBxeAH7wizo4Q1lop+A7NqN0O+RyndytSzmqDRIfGYpNeaRSzh9TFGOJ1
4QVo6CNs59NXmuOMmnHYB0TmgsyVFpC5zNjEobNA0e5LYARLVcTNsbU0OuNGwsmZlUJBQKLyrszh
wi6Bozmp8KhSRQbxl+GmUIRMIxO/WWD5LclPyQnKQ+JqVEqghtK85H1poFbEt9N1gAm0hChP3dAZ
y/2Qmqs2OMp6Xxya2kfiu2pkucvkg+GgzhN9OMcpspbgNo/D1kDH2nzpaa4XA0n/YYi5PvVZatip
rYrWrQl6kkAnlVtTdFMZfknwCCNt4GOErRrFnAW1H8qeWF1VFedtP0qxEhJ3o33JcWutM84a7bNV
hAK9mk6u2WBe6Y3l57xWqbVmkvMflw2+RUy6rvToCm8Nd/ijfakQYJMoqKztMuElOt0gVaddCeNT
nvs8CXXi1M+EPVjlO1oz+Mj/BO2Nh7X5RbqQgKL/OgRbm790AQE9UCzAjQp9qs4LBYK4Mc0QUN9z
MqADzVvRG/B1+QLp9cjIladUVCh1wRx6pVhl5T5Uwv/dJmw+sAWwYQ3fdoHP1omZsbVYO87Prga9
LM1/qDtosuE+Omhg45Z7gRGH/ByRqb7WzIKV6UtRigvUSYICquTBwlGxNaPxPOySX41PDF/3Ko0q
IovGsUu1/gKFI5RdtfoTK63bF6YJjtLppIcA28yfcRjUKCnG4aBAqgVLEof/68kdSPe6lkvKoC12
905bjXRUIkswRZ6nOoFKWSbR+oJng6Ev+nPLpEndXcXacc4r6k7t10wtMh4ky/W3DzPVE+OegWgm
xRK0Ki+GfuuRqgE7PIIGltxG6YMbYT20tN9SbnicucGWszj0l4uyjrgJtknFATtBuosaJBmrMc1P
Orv/Kq2XiTG260qlZ4nrFDkN4HTDmrZGDUtOPxvJpeILXRRL6/7n8Qnw3zUPJYmKz12AkbPLm18z
pj+DeS8T1ggZFF7zgald7ElTiL07CNm0ptuw0Mdx2Pzh9JKrz+y/dAboesfykvw7O0V9kjuy1JZ4
Aie0ut4ZQwdMkA1fNuKmagl8ca9sAXn7vmFwb6iPDQxMxYiXlVEuYxBxgxt/GkcNf3YbeHwcZLJH
itLRzKDZsvi9NQy/updMKmNTPa1+u672UWe58Q+v+SXOBCk3cjbGhJsUp/fAux4Rac9j6CDeh8cC
UbO+9F7HR7yDreEUXoU6TFnIqIUN5qQkVGOaUacueTyK1YPxdOeApIILJNjBak5OxPUJOgeDLwy/
s4qR6jd3e4k/2Ny6HPVo0iltykkUiXpQY3zrECLWgm7YsQPflXxVi4auLV7lw3WoF+/rlgjaT6pi
Mp29zBmN7/Wj4WiktinPjkw8tk6MroVjHlegeuGjvvd6O3R5/2eUzJtFquzRbILJiqshtm2buGvt
7e1oPLj4F/0SMTShYk6pfMW9DaA0uj/1MOhOEHcnb/wSpBJ2xOTwi1HLJ3l1ah4RV1gvdj/AAimj
T5sRCKTG6Q4qJPK1kYAwaH7pyZ/fi8vHMhI7uYLsKS2op5KAXJE+7tP70lSJKDxut1PzfpEkOtH1
0c/alSW+OHEgzaFpE9Z75t1c11gPVJf4RYFPT6KFd7Mt/aeuIH5Zzzv9y9H8LWPWFGDFj+kACKpf
TGXg0VTfd6UKPAuETVB21Oy+MgtnoPvv83Rnfaaht34xL5TvAyMz7W0gsWHJxLuyNEEaCSDGPHX9
hdRVrA+3ObTd3R+uykyZtYYGTq8vBtpPza4CiT/ZrCV3ZG1wTd5WGprCJjGVvlpS4caVrHtvUmj9
ZbmF/kX4NXr8eRnzsFGvd1wo6QK42xLJ1QAUErHg+DCNbYzxg/jG4DBRZNchhX2RbvRkTbHceHcZ
jZYniVepF1abNfFDt6C2D5XIFV/YkozSL//0AqWOZry+aoiEQlte5rm6OkaP5/E39YVWYNdap5l+
oE+TaW8444HdSNbfLpAEVx2g0Ez+rPOXyWTTlfDpU4rST1F5Dcv/hf/2dFD0Qth5MKeMM839/xQh
5aLu5Vsnucf/5UDdZqohHwglDUl8WQL4AoLxSAKLwt8GQn8jGJJ74LsQ2Bapgtc9rCxPWNjYzxV+
AWNrtZj/XrOxi2GdlqRVCJekwgYjWVpBy2Z1bf2/BYtL8djuOEYNN64qk0p8OpLxXkR4fnL2S5NR
w3FZsWx1fKymKxKKSZgikXdgosJzi8aU7raWvRGv13c3AGZMF/nS0/M+tsNHq3ojhjocuV/N0WFH
Z0X6O+VYTrlsRFk24yDFY44MiBvZHWG/giCPDP2PHlE5J0VMyaLTQtA4itua5F3q65BZ0Y/hKz//
fa9XQyerCIhMxQV9vX7BGoG/EKuk0VuMwLs2OO3MvayUEF1uX1WWNATCtEg5oNLXR4ydTsR3lYJb
4NEqonrJZuno8OEKTXpHti8BDSHT6tsUtIoT1hmevPPwYkALuReV8G9+01rkJLR3YFMOFDfinnVP
4Y87CeuH60GvYmgonMgIHysn9gCGuQwWilEW4sse7UcNbtO02L4OVBh7FdDlvThMRdqreBsxN25r
Q85cw9McuhiXizGB81kjjnAVS/nEU+cHOBSuUFj8ImAICkWajjPXZ4FVlHaE5zki7iyUWhyDxYxa
3p2eDDsp95w07lJe7gAoRTT3qvepVLClj6wamm/1fM1VqND6sWwPI4G8F4l66LTfotCgVgueI2qH
qcqr1UgKzRArCqGDM9ptduYuZIkk7zqQPs6MCQ7Ogr/NtDpWTOlcC5neo3guNmjDHOer8T6rUV10
yLfWJHAjDa4P8fzpC0x3HP+hai63JegjhHm1umBuuwy8kyatB9o4FjKKI6LBqQycso4Egm7vYJGw
t0ndHolJy0MBF1/t3n89+GyqLHpxWIfzciE6uyV7++Io1h+xCKOKPQLoi3G8e7RpMJ9+2Pq4neiy
0EAHVIloDqXfkESHVa6lQrjnuy/vNseZzXbsJ2hZXZAJeB0eRO72OHqNI8DIgSdRJAIm77aeyJQw
1Ol2DaEOkIUm/J992lmRobqBk9QNuBT0fzociX5V5veDwN14P5hNsPWNeitl1ebjxKZjhdusK1lv
v7pf/QtunUv6jYA7md9OdkMsbIHYC6n1fI68MSkHgbdyOVHgesrpKfXgf/q/u1ULtd/PVUnaYiG8
k43JCJMsmzXlEWPttVmHMwfXScBDPsGq7hMCtbTJHtaydprEhuO31snxjody1eeYUS8fPQz7OdVY
9z5O0RtZAltMSPQnv2AH16dI136vBwmYoA56kMGe9uqDgxSg+/BXGzd1xVuAVXGiGv5F/EC44Ann
KMS6e7LCIeEQZo9PWKTRPNGK80IVj0JHllfNmDzolkTisj0y+oYYN9AvVYfZXaSp/n7nwS2Cdpd9
qDyy9Pmcpwqet0TT7Kg4kElmV9TSngsUkoMW8bV03C+q+Peh+NrXrXOfL/HgNg8D0j4vG5T8HTOd
J9FhLxUiGm6TRVvgdXu9UwfHQdK1zMpejZM84u3UY1TfzUqXEc1ZvadbDXVpr8fgJF2Pb/CuNcq8
CyuDe91ilouW3ogZDaHBZJrEVjpepbYTWzrt8mcAhQz45jZpaImSToFoSm2NGmyDrsQ6dbB2eUy7
51jRWkAGv4wEZkolw5GhsnwXys49RK4ZWMU4INzWfwVH6iryaADdaiRsPCpIGjgwA+yc6LdE2moY
Q7Q12Du38jco+ptHJETOObIu9w4xdndHhy4LtpIc+0bwCj/792Kf4CknuwU7nEy2ZzPsAeIzrU9o
n21qZFRVgSI9JVGx1UV9nTJ+1xXz+g+8Lu2xT2vKRdHR481UinVr855MW++42DS+PpJBJiDCcJEW
RX5O201vkg3wavsi3RZc6A9x9N67XIUTJCCTZ1z7FqnTzjdEcGZdcevEaf47nqUAWi6Fpv0nTCzK
vykdv9HmG+6QjOsgz2wTMtSLQWpOGKOg2QCu3cLczzjRld4Pd4QHVpateivOjVTPUfc+vgc0Dnh7
CO28ySdZRFItiTqLPN0G2nv4aFdGDDU36bQw4KD6FiB/Ce6b/GxQfS4MLSTdpCtbIQIg4R0LxTUz
kdf90XhdN4c4M6IsbpprVM5jvOZzHvIbWa/kxKqgWPyl42gRdtLqedbBofs+BjgTXlolrenbffC/
0LuFBK0YfQ8Plkmi5BhDAYFwBfXodP/CYfUn+R2Y+s/DPxM7FymPJAR7iNoOvheIxdhLjbDw3S6u
FwX3t9KmHLiIE711vlKL7gSTK0Y6EaZ76pXxcPPIRKAMuew0BZPNUjEpxtDfabBokk8pRUbtFnzQ
x1HZebZYR+qz53ZrRl7G9O9KJiOd7mbOzFeF7vTCkyRoHQzHZjccnZzjALG3xMfaRsiPvinvVgfW
XRHJObMUBVaxfXQLXMDnEWgGgxYkQmTOshy6gLdEDNPySJy8WyZJDRTcmIXZAPjwu6V84Koxcl3v
gAykLlH1geNH4PUrwYldkxJW0BWQEIiOQtIQaocURMAseAjmhBRc9djVVJFbNQsq11Q8V+/MvlPV
js+ND3HBVMqy+3u1MN0HCTtKEYXuSm6bhsaB7UoK2/DqGBjafDkMJ92aDVU1n7IFWeexHA4xnjvb
W4mGEo1CAan3DLjt03dDDtyCflA8ei+UqeqZubL15RJEL6kx92pVtlY9gIkZ947NVsF9nGYUk3iB
OqmNm7iJW2j/lEvYie9/zKo5mZxpnIv2YzFcPcE7r8uLcYO4am6/TrUawPg0mw7NCZYOn799ad/n
FMg2g1fWJzYa+y3lJPDPkqEm8W58lRRJTnH9Ll5Isy0mN6IoHyrz3iatl16ord9zTU2J2JiNLiQK
W/Fo92NeT6HjxMLHmUk8dp4S/qZk64XAweTxAS5eHGk1lD+3wU1g8I708R6lw1hRnB3xCeBy14/Q
nlGrD1F407K9Lbo22qNEEMeNUQnQ2ZfTS+0nl+XVGIfFB5UoKkAI66ya5PfMoJjkJ2XKT4IUWJEZ
zGM0cLp+vUigac1sP9KQlQ7wiYCkYG5KEhSugGEFQhvEx+6SQPPGXir3SJvl7ng5UJEAiYvHzy2A
XKyLpyxBTeJf8wl9lC2BQcgd5/PjzfQAqbKZigQHbfMC+prS5d1SI5cbD74rmFJ26UAYuzjGWQvk
2N9JM8wUNQomhgM/enMcwZS0r8pqWET72EL9Ux30gFbb6aqbLaGndS0ymcjGlvA545OgZbJUSHmo
BDYZ10T+NXTrT+slRhbrAHCCaov+6Tc7F5jQk7NxRhdqi8mUi1WBB5fXax74xK+tFCH3EmGr0POI
AF/Vdwep+eahTIxgl9qy+xleGK5NFLGfvYSNMtYv4qxB1MWXVuqP92lVssE773JhHXnHRI3zv9/I
J27UVRXsxLohniyJKIFc2WD9YauJcrr6TCs/4gIlZb+KINpgWF0Vowb5mxDwyEC8/P7Pjp8CjBMT
EzxZjwBUmDZR+JbY6ax+urcpieIAknO8JoWtBL2NXvKM9qFbfjh80EeD7FLbH8WK1uKYIUoXKiLU
5+uSKnn8kjz9TLutRd9DyoDyllaTCtsIj46nPc+F1sQRsULi+Xp8+AAZBpJgT/qCgTuTbLfvmCeQ
V+1WYcOiWwL6+5CxD2nJ9SKW46+og2ManIkZCZirNv52mQnVLfh5tBUzrwXihKKl7E3Xrx1zSJZN
23lkl0G1tYksxToliAjDFEayu24z6f9bbCIaXXo6c5XdN/V7iDzzGRKFXMqMcGpJpe1QLR8d5yZ+
R++igMkR5hRMLjvtulbIVFJdfsujUSSf4JSX8FSPiKnXBY0WJZtA7eKrrd/mYyP7bJjandQTRPAs
5Db/4UighrhjrRXr98r72BPMpZaCGTa5S0xDJdHKyoPl31JBv0DOgwBAjNGRGyU5FZm8JiRu94Ny
3gUmKTK3F4AxpUK1iTaMjmFYWdTCkiVqQEeOKNRs3Ge37K4QsEW8p75th5XBe+ejBAcNa+I0CiUX
axwrtAM1Tq7QjfeZA53hLs3imHezQjZJ6VpFE3uSMqA1TdSk4E+qrw24drnG5c9xAeT9E6judAQL
qx0oHpDlPPyJ4TdrAPiqY73gUa6qC/GEmZxW7YxRbPByMcSDY14bglG5yuPT1jSePkxV0ChP7jzS
5V7lzd9kRP6RvYpxlaDajDOHUSZ+AhHhi9IefhfMg4N2KBRrKzV4JLIqiV6SG+ruJ+X2CH3zPJ9s
r/Vp7u/6u9DfgwlJCXJmY4PIVBkUnJCleE9/YI3ytMYk2Wh1f4cnZq81CFmiSGH/86mSaMAmT3oC
oxVZysuUEWVm7GAj6v8S19YSz9y2bCh2v9C6ofWlOOT6HCRTxY9Coc1kX7zxvbTDYBJuQvFVB0pR
gwIhO7mBCNmY2clN/N15hPCUyKDyBuwwOdY33Zq97H0Gwfu/k6mGikRYHo4vslrK8WPZqQ5gghRa
EjngCWDMvH9n1sGmBY5e9jrvNt2Hk0VQzjPn2ldZZlXcwfX6l8AIO7Kv57EW+xsMylY91hp4AhDs
8GhjuHBDEMbj656HQ5o5J8AsbO40JRw9a6hw/FWGlqR/HMXHdig2/XfrzIHrvfv7niBXGNNpXbl5
ZXYVA1LgVE4T3Wh1Qs34Nx5MPVlBUebq/FOTr8CZmZFclTVJGZ9V1tjDrOFTqAvRG8eH2jpCY4r1
mU2hjUm5D9OOZZsnAwWgGY2AK8EsfMkiCLmNSKfUUAPPlXL+SmNGJKAoSNfvP7YpqIQ/n6tisDxi
MbNExjtKY/o3z9WTbuxX6nEtNyPm+Vu/gAfIHpyFY4EBYv6y0RGuLKs0YYi1mm84AW47ZA8WZ8+c
dVNAfjsTjuvOuRaMBrZ+2CSU0KFWcGB7nspUSV2s1yy7VOEjogjZYUgpXzXopdDf+aitOs1i0nqe
C+ehEcxAtKHrU15wZy3AKmvPIX0dh6Pd3W4ZInGHdTCrj3Jqmwm0TcQvarWvLnhfds0cq1ezv5jy
5Xv7uuDunzxfTZfWWTQbEvPq+CSxAwH5HtRd1ugZP7MAfjH63v7TbAf1sS+xWdt6HloLiObv8PAz
6dsMcPc048ev3EVlIgyqG91qdTjbiq/weWpWJvg2eZQeSZOkDwfvRGHjnh0+ZzAi1cl+XDxGhGLp
ad95QyR+xZRZQlHGXdwlgNJDdXszZeDP/1oZSGwSFXIjvFCF5ku1uUaPua9oYckqEm7EwzoIM2oN
ppKE8lfTcywZyGO8uWu+k67cJs8cw0nySnhfHacFSDCjwCSAIvZhaDoXHVKeCWDNVBP8gXX5gZip
p4joC+FgbC3PUGphvB1H35zEYo+pBqr1w7WA/JgEEHqXnMeA+55avI+a2wCC+tGFlmsZfWP6l3i+
REIoJyoiZb+5SVuGiVo7oAHtpm9UXduvXhhykSbbDohBwJ7dbv+kcLUtHouUfm4K97mXr19D5h5H
/FNeMhZJtMfEGsHtFZ1gWFcvXtJyl1tygWzklJpuA9XhK3NlwJ/+fLcVozuFpv2YJb0P1GOAzMk3
0zDoPDW6uaPdVoNdxI4ONEfFNkrsEdndx1S8K5Hh08OOoteLfd3Y/v3ARALeMZMz0pQ+P6Aujkfm
q3E8GBz5VILR9a7L1lc4W6BZELb89j1UDxGKrsYyt4kwbqx4A2BV1RxmV8lWG0YlBWZaNtwZGlcR
t9k/5loTuOsj0ejUucmy9mEd17V1VeTBaJ4yCjLTGDdBcpw8nTgQv4fNC6NHVvjpaFWdgL0A+U5e
1Md3nJzaNYg14rB6Pdttakl1H44CPF7yD8mL4xDbWeznJ8wyyTgKKOHgR6ApX/tgqa60JXk702KS
0g+CuGTvDUTR1uboIRLdYR258bJFBVlzGAg0pLIeW3hRcEf9y9G0zWGnN44eCDq65HARJ5QAe5mz
jGICaiqCFp2zi9PF2Vprgl0+RUEsXaqkvHxaqHVRCg1ICQd1iwVO3Vx/FbW8GdMDpq2vPp+1ElMg
sdOV81YYtWGysoWkAASI77z94/2B3mgpvwQ3gQL7W0Ajy/WcAe+lc2woQmWZiGdrNwBWblMIF6ic
dX9+gVmbm3Le4RxZiBNAQfPNiYhY0RjTw5SuojAjkngzShdPq5nQqvjHohy5/lc/6tu0q3qDl3Z5
oI7W0YDjrEyerogS67nYszKCKgGay6I3X95zMzZ3wqf0PK/wofI4aAP/7JPXK6lIE29tfsjpVSyS
ijvWcd6ctx3TDd6KuJ7A2ih7nWwIWYGgtNDXz3j72XgS3MBRzFFmL5G377XY+0q9iYYrKIQfRgyv
oZusZBR0H4/TcVw1NXP5XWVkSrxgX80Dj/vJ7g6Fzp46oxZHS1SWx+8L48asPgpP0BArdd+VM38A
V9QGU3qPHY1i2tsIYhFyzKQRWfVIVaGAr7vvq767ZYR2pjgbQ20Qc+LePEyMylGmoJ0I8PRs4jSY
5aRMUzeg3GkkBeOIZ1Cgzb6KUJUsV52dRIsLX6GNWw1cHFFPz1dpmT9OlmptnFBST946El9TJA7x
9mSYURjsxzrA1taEeRZ8vMQw4GzgqXuQDKm79yXfB3AxvdHPY9DFGnWe1gzX5fiWhJv6QCSkLjRE
N5SkHIWJZTA7eOvr/YafJ59w3gAbXEsmjoIzqC3vUcStdTq1I5mRFL6K1DF1QwuJq0knWE2au4q0
PQSdf/K77LhdhpbJT4w6byTkv0iEH7M0dHJ/LNPkxWelkJlD2l2VcrTvbRPbHHUYL6WoENms8p05
0iUnmjex2APbrL/wkH/C7Knh3WuqCcjuwbai8nwkDAnzJtmuZgSayo4LmU9FbPNm/ycosMdP7c/d
LkuRThDFILtB/M8JbROM+5h4yP5dhonMgu+//rcBf/nltpRIfSvxG3g1Jyvdc61Is3leZON2rUSz
Ay9hSzS4CKVpcW9FxdxNHwiQ/a/xCSR5k+GwmFM+RZziaX/dOL83pR06G/oB/eW3utMPRX2W1WNu
5yR01gQHp7JDCWP7Rz0/7y/+XbVCi4zSw5/cTK+ywHTEYwhJ23/WDEOIcpnrXrX0fyNH2KMAjn+R
tGm6FnUeJbw+ZO/nDRie/kyK85jZl1fpox2fcfVVZIaS7eLZxFRs6/WBDrc+m1IAYFRSqzjP/ti1
I6Ne+sPF16aVvB5H1fQu79Nc/cn4B8BbOVywtw4ZWlxpMy27a6cPN2EE6GIYAQGLf/gPUAu5vnv0
uxnDdTdI+efyejcprAR2tANL+yw4q0N8MAIp1Dofgiev31kIrRJ1+AqdUQjUqsAQkFbTviTXArNF
tvD23iSfJ1ne860udr4kAOs08Kk2jcbNJp2SI9akhOwBv3Z73ZQ1TbzW4Xk75SW8VrcOEFQxrENG
YxtSWBl/Vhky6GRTw5RKeKOM/81TMQcQJYLsHYk6gBih2eSYo2IPR9cjmGofUd36/H0X/YNp98f4
jnYUYYk0rMRGVm4rDPTCWeF++E1p4auGEu0bJ8uWAM18cdloWkGFn8o+cfIVEQHzihli0vc8nQRh
dlyzZZQuc//EIGaBG/g4mg2bxTi+hB/ZEU75vgCbyOfL329O3M+Iv5SCa4yMCqUBxPpbO4T+OD52
wbcR92CuJ+TtupTpySHJeh3cHbyZq/F9cJglSRZdvkuxOYIOARDXEo3eqOZIDJbiyrLXmVUDpvJ1
F6mAThdQmRO9U/BE+w5p+Gym8d/Lp42+3HDnGh/PpIQoYB8WTFicVp03J/1cfbxAcTKh39TdT5/3
L0QphNU8Da4ZcY6xMa53TbYeM+SNbyHnrOwv14cC+HRVnZyMI9e6aq49uSU3m+/sXpxxnT/FTaOy
xDVSTEhhZfVV8zs+9HA1Tv4BfypY8mI3U5MBBt3gZAQCj/rbwTajYk5KwjS/RFKVSsJuRMiDu99j
IgMOjXRx70Z68UFaV3iyr5JbeE2mYl1HwCvMlT1wmW+cws3hw2ZD7WIP0NFPVargaIp1LMis/0Je
e1THPUbZPc9XX9If/0FIaYXg6m5GqOH35fWAAnjMTFrkeGOOc4iK3bp6Gbtvv7yPrnt2uBLndQb1
5DGRb2zGdE0AUK4288J74e79bndI3krLYAK8nOZhULzjYr6e+twt7PktBHApNSSpbYm0inY5/6XO
2hvhjNJ63Xjwk+b94lkvNhpKeDf9jPeHFgfrNqh0ec+vU0i08r3tkJdJPj41XCsMHms4fHEEdv44
ZcsJ0w8cPfuLCuDeS3fuv9j28Qf30Tcvl/DWSm7j2wsSueR6F0lbblcFyVopO/kczwASNCZ22zg7
k9X0dS+45vabAuZFoAzGJLQB7O+4nV8bjfQUAVJ9D6ieySr+fJ4v37bEgd7kg6l1qVJAgpU3mgYF
1iweWYiTcEZvSe2nA8oPLxZeFDWKiRELVlO3GaaDsEakC9O+VsUTyxoPccfsnOB9YD3wVUSzl3RB
9kqSR7tDfYc92Xzw+0q4JmH3SJEqpujsh5iSY4NyBFCEYbWqe2ek2lEJYE2xzs59ZjgV5OfKOosp
samlf5BL64uuR6iizuY57v/MMPk5WDPpoKuORsnjrlNGc4SjszcokZko3d38axC42MtkDYjWrMVg
MQQ5Ff/LHLrGdl+6IDnj2tfqS/RNCJmpBKqsyBjYScs8AO915QtoEt9UjWhk666KXN9v50gFiMSt
s6I4P63pv+i1kIujgkn96NOM+NEQhlGWRCfzGdSKKuJeen1q5JBH6+Z95davfZYGFo911Z6HIgGp
snODaRw+FsG53lqOCiWUbTQ2DvCaHbT7EydVZdmHRA4xUlUoAi343iV+BTEbojOsApUmK1BmMIy4
Sj1pf+VuBvUtCq6XnE21SUL7qv4jN/nFGre6a8K2ZZMZl2Y6IjzNCphnXuOcaWeqHiQU/SRNDi3C
Ir74DzETra6oyeTMqPkq1W+fjOM0xuI1rwOkGQwUMLyyVfGC8NCZmN0o3bhEpUpKluMbQqxiDMhR
Po+KeS2FvMxnjXEuBkzgB9SJ3GEKm3Hm27bDLQ+BVCYSwHl6uwowBJ4BF/WSyhSHGQPizssH5MbZ
WudzctTN9l3VJGsVSflAoPn7eLY9ojGxf2eJnGbS3ldX5NQdFRQ85DThuf5hdBIl5UScE3De/pFK
amGE37GUd1ODVPrgffqYw+Y+YLnD+rhxStthiUlwr5WnLHG924CmIZF8BF3TlFn16YHUZfPEmlW4
sZw1UjjyBj+SQnMBIB4dq2pI46829zXnagQwHshubDkHbftYrFIzQGVw4q/sBuHkJBPhGJg3ekkh
tQXCgmid3M4i68c7FIFvOwYh/4Lt9aGy0K8lE4huf7lFlTlgimfJTG0+k02n8SRmB7Wmo4SLFesH
qxueVZe/3wJYyMiSfGdKY2tDQBU911KzQAg+ePvxGFEDSBCt0mWVR/htGPWbW4tQvAhjJIYGFrcq
9bxsG1qzCq8G4yO081m6P8rEMerOVScXRT6H8zyP163HPZih4XNYAmi7YfwsULjo5wdjbuLAs9LJ
TlTlv8ftsY3hQ6OMXiS0nkzcGwQS70aADKdgjruP4sgfZgqnp9PxABntdmM6gNVhQHrpkxs6Cb92
ma8c5FK4092gphtiIWKJFS2ODx9gVITW/feRiJqYcx7NZPddfq6kbd9jJcDETqvieJfEClU9H5ho
qyQZe//LJtkMD003aU2pONLBnM1pLboHEs+2rZs9NbWil3BK1UZVPB8LN1KJ5aVAZ+1cMzGzFjyB
4AqmAsL9MAFv/xLSqqdILAE5mkMcRXwagPoTY2k18fRnEqo8hc0kw4k7ZMS4AJ+JOvu0ijaSq1I+
WnzT9hzqrXg3SQznslLVK61OQiouFE6B8y18zlQlIOTDUZ3mJqCO7f3rc680EaxnA0w++Uq0//zc
RWxFf+RMZNDbfwk2timJgWSIOMGIpLTErYlhiK79k73M4FOReauqcNGLlzBwhyXMsMRZy4y7+rgs
HlZ54bIW6IXVLge6HK9g3yuBA4sJ3tq0TODF9Hiy0dRo5V5ST8t95LsePn8oaKSNRXUEyKM/QoVx
RRiFbSilUhSe5q7b5MWcRnvjz1ggdY6DdqyJoe31ns+DBQ7OD2h9FrUD5FG0sfoekOk5ZF9xCoHn
uucObRVfmDNG/45tIrzROyO635om1LiEHByX1oBXOqtEul1gUeHQZcnZ87zzq5UyMWid+upmJOdY
+y2b2ybyLrq6uIlAxWuS96BHSgTdo9+lSNqP/sSxccMtdKSj3m0sI0nflaWsFo6rj3M25vNpfcKs
FCAZJYDxaAfGhD6J0WGippvawt85XS7hN/no7PVDVoYfxLYjS18pyp3RX2mVmySsa9DqThEdSNRe
IHyor/AbPB4XrnUW8B7MuMEb1hsbp81jfmhlVnGWOgnitRIADBbhT5At0sXdX4QvaBzwrjgh193P
2eepyj4/1R5lwTMb1PVnTd97ZGkY/yMdDXweKKkWFF7+QFroQ0CTVp2JW9n5hIvXvbhQL0U/Gyab
mSvqzfN/7W4x+0FBLpfVTo2/jEjJAsZ82Qzxf69Hnr3wwxW5JgrneCmViJwrwrgScFKe2B7BaIhH
idybtAqNG4HlxX+fvw5d3GSkmSaJAvfSFm3fbU1xnqE8yHmQYZqh3DwxTGGFkZs7aju1afXxCEGy
YCT6oz+lhKW9Wd9bZrzC6fSJD3OJsRBzl3hNmjC+2lc/3d8MY346+bkZzOmf9p3QD0bmPL3iWwOI
4qmhUDfukJhZsS4FJZfZicVc+eq3u/AoZkKz6CrTAHiVCYyoU4xvKFEpBToLDf5xzf6sxQcsmP7F
jJU86qlj6hupEJ1z7R8lAYomQiAIYo8IkPU0K9pkBA43TdaUT0Kc79r4QosUVV36cQSsZg8OhWgj
CfE/PmbtAkjuaGqq/TR/T8M1DApO/S585Rl/Lc1P+kSmzNy1yRQeJ9IkbgandhoGGVUUR9WE1xDi
c3g6qF8ryB6jumYPkhqlNAZdRJUVx8qvAzSVC79I5eKbrtulB5ZbGHW8TJ9+RDliD3O5w+5OzSbl
eSYKBXcgP1M4AiIB8q0CEvmXSM44USUwkxGweza1n0GeTBx73+WaekKaI6t09DMhcgzc8G8YR28C
lpz2pf8pSdKmFIGui0vcRzYGRE7QHt6yJed9bm4/SGrmpVjez6VHTvkzq3v38YXnnmKQ8FU1KpbV
77pCcrd/rje6rjCCC5NXmIxORNaj01uMFagQzHFpW4dKLelTM10TWlrL6QvjEaPswK1bgQ9L+/CT
OPDiDeekDYf2uLfitcrd0aS48UsgnbfbWoD6W3oieMW7DNsPym+SD1ArA22biE3MYqQJue757QrM
noQJXcmIOiozg6yrF2Ga3myA6AOjh3W24CBb8fgqYHZxh4vamkqkzarJxGTXNg8HAPV+JPlaVOSs
lEVCEtme9x0IATWIdp7eYg1xhzanuJx9e8u+GLLlhMeW6kdUbxGKhb6P37xofeCvfXh11QCwYHj7
BAXCuoT0JuxkIT1FtyNKNcou/DRQ07RFnldb+nLTUNOr5be5qxxTtUoXj3dRbCMmmQQq15s1ACzs
rnbQEI/GVcYPct2fZaUvdBzPgVpCnA+9Ra6t+HwH0daXS3T5scuBbeI7yWKwlEMS1OnOm/5yRtpO
Cp/lVY7zy+d3tts1DD7WIqiyyWvX2hYm7VwHVYyY/EGjPw6hhW9nRt9/GYApjNCPrW5OItL7MV2i
WtjWDf0dBxGH93diUIG4Ik4hP47iW1sr9VxxrAKdYsYAwyume5somphZdhvBFCQ8LN8SE3dLCJyE
i5qRXcEGotVB/QYGDLtB53J12PkKbuqM9Hm/hdg+0EOSS7lqCN44d/6f3A2e5HyXnI98eH0R6AmW
mtHVbDfJg2NOk0fyBwcg9llpZJqY4gqJTY24F9vAtH6m7ppc1Vv28flfMQ/B8eKeUx79hcVN0s09
oX3VBQRmTY/GeSEIjIISM4SN//iVr6drqaiHsy3w+kZQS28jzuekadY38mVLvL6TzyP3C8yz+rLo
3F51+izzpmwpJJFbMYXL0M2SMsG1cK9KFf3kLvL+ly2PDn9ljaehlodriP52gZTZErarKH1VCXaH
T27K76rBkdfuzEopO62TRQdLC1Z9/fIMoqp0b+YLV8JDsLzdzLtAm6iJzyNhIj2eeUDCiZfMeOBj
8DfwZr7QIPw77m8z1/uXrOYyrfprWW8Jb7N6rE0GUGK30sASoClRn36vtU2G6IIVctIaX7/LFCyz
UjVaxEVKEIHmMRCwKth8tdDX5PUDcHotvGT3vJQRztmFzTBZjL6Rl2smcHmzg/DAsXBv1d8T6TVU
Tm18hRfgJFAmRc4q2Ol9BldtOfB++8P947+qFUVLsL6NVN37J8SDQOgiXdrhCOqoLkkUyWI77vg6
Gw577IGbs3w5AP87f7KwkymXpU/CSHqfp2rxzPiGv0DN6acyEYRND9IBmJnlBHXjk+CxUVka8vtG
HcqpGbOCXQvRTmSiT+oIi/B0zQwv3/R/I1jyp45W8gLD3KO4/oD5smi8h/qFf+/PjjD+lSiSmpdf
Fr24WnnE/G/SEiyLxqKc2Yl/5bklsT0PPy6Zdx8EcnXrMZg1/JCDzpe4z+FmxA1UxDl26HwxYvy4
CF5lRjxSShKJM96zotuNLsfPRznTUoN6W4W1RRVYaokX4jti1PKQUAXGvFnIKR2n+5Dfk701a3jQ
FjOaNqqDv2edYo1hq7gHmeuJnu/bbyJ6biY4vFjVtfdVyEbS3GCBkw295MaqQe6+L8C/F7ckvd9B
we7XQuNHUDzwOMPf9vEukupjzg9FovseMFTnhK9joVqGesyw/szcDj9XDPtFFEks3uk6od+RbBWE
zAMdyD0G3T+6d/QJBakPFxAY2H2VGVxiYllXzn3YhZnNNqdVTMvUcmxqKt7y0Efy1oQQp1qzqKdA
LJ6SSUFHYx/cwNPgSaukrxdWbjaPFQD5V01bJJV0ieEMa3R0HwUs8zt9cKEgk0eUOCtRCNEYXKEd
rpKfB7Jvj4vb0U0QbOR+hfQzeUbmw3zELXHgV+yPaqPeIICYAyMDqR/cluA3gM5Rqp6vgTPMX4II
Zngj/xjecwJxU5Xsz70Svw1jC6cmvNtDo1gi5AZQptzQSa48R8n9H6VNqgv6r4Q5t8m1HpO4zphw
vsrDtUunos3q9cga6wiDtxggj2+a6JOyN+x1TjH6wtUcipatmZ1WMs4BzCAZQs0kOIYC7Dg7i3cB
E/9lfJ2EVB6CWEAnYK2XJE37PS5UKMLXTpwQf6yPaWTByU66UYMygKgfC4uzoEaYH582CQDgF/Ox
1qCRU4Wm1W/PAdglTsJzQyV8Rj9h9e3NdS8V31H1x9Z38OgE8hja/aGoWZLjnXcd6PkspOTJOIip
ARvpqtkrxypuPcxJy1SLQ8ykrfBfkRQ4yDb1mkdryBA9RsnVvIV6deh6wDCjhC3HQK9HEYkKygEM
GaeMBvh8maW37pFZSZ+QwmuktB1CxU8Mz4DykiPe4N9WFP4ljNTAu1YJgn3+tq4JHvIE0D3YbCcj
DooKdNkZS7E4yPh+dNN7wYfWlm3ZBnilm4A29OHNuSGv+1nJ9CgxYmYUmK6UMeuht+np5hBtOp+h
WPDsoDyC6acs8Sq79y0A95fbgvmIw3G/d1eqW2ofyrqw8sR0Lt9TncAxRnLKinkycbcoaGwWBGp3
yfmvIYwZ2A6N4mE+EV6wmitQCKTBDHqdxsfyDNC7adQB1dl781IZ38B4P0Gv9fI43K/+RB4e0q2o
YZ/ZMoyeFGLr94E6pqoC+WuDjoBsFg3t/dq2+i/md47LjPgJfVy9myE0x35osCb30zwxR/oKYt8P
EtohEQXWa0jYsx5KbhJC+fkL02Qx+2xVyHOcph5xBKyCEyEJ+WAhl1XoUmsJDOTrjy1CUGIhX7eI
SjX5zQ3nisVvREGMQZ1gGn+u8KsbHcEN+bKbCbr+ZntvcYnHLV6CkHjfajL4qpGuM+nrKndLMvAw
+8bzJiUzFveFsSc2/W0+ZguXlgNBG6PzcniNBpeAjPNIMJ6sZAV5sD2BAwKrJHxvX1FvCKsqTbPT
y8gHRNZvyUrViTLNKeijPCzU5ZHjDmuRg2T/C/t2ioIoYvYkfEWCAoe9sEEl5wvWOcmr1orTkqh4
hIcIPnmBf/ti2sf4b3TVyaJpWGfoNpodWnrHI5bcJs4htLKekOxs8/wTBFeu/JqaV1Nwu6a+LOr7
Hb1586nvuVY+4SgGHqJOU3RFAcmNBLbi3ohzjiwpP9UgRXxTsvr3SNu7750ntSJeQX8Ts2fz3eJx
c4PWvO0UVjJgjUDFXLJacgYAxfTqKeyTe9/avwY4hCJnojuHgYjtVw30mb3Nhm2z+TOfEJQrW3b1
LVhuRcuFlCB5Srz61Yd4iUNOUc2kS8eIJiw/cIJPG6UCiNzV6rdHZchb0q2gAWWo0PqEbHyM6u6W
oJM3XVIVkm4gJ1tq4XqRYEPekyQX2oPkmt+zMIIvsKMlH9A7ourCeAwSXifpQk6bBKQQF4kh444c
yz9U4MTPgL2Om7DMsxlkNFpdfoCmXcH+y5pOsUvK5C8Geycd5oJhaf/9V7SVzCYQ3WMIq6voVa7t
pbsTzOTdmpDfldTsyyIoh68mxgxhDqYe14ZGfyYjYD2gIcslNhOR1n925UNArG6H0aVDx6qZrdCq
GFjOTdytv3CxU0Z2QL504E7RuV87tNaB4AFVqiY5Xz8tJD10R/kAC8CYz+vjtPjklQrXvDXSipfz
cnIX6O2JPPtk1AmufH2Is47vNqfCinQoAr25kGmoBw/nGRHFhJmWDbxQdhqjShSahgdtaSU9MdF0
Dj2eq7TLhnw4wHsOut9cH4gxbuQJAo0hjAG/NPMFtRSN29Ab07MfaeXiu+eaVnXPs2nC92obrPUd
0Frki7DIlSt3hWnTzLjjn7YUH92xkRdcjICv6in9NIYNwXqr9SeiDALhJMZCfcnKYTNLII6lQDOJ
zJmSshsTNQXwj+SRqCIR+WUJJ+2EXiGgmqcC0vJ3+MTXVI3hygL5S7LFRWNXPQS20LADzxUOIyK5
4NguoALkAZUG31m89j3p+85VGqK3iUf8CMkbbVdsiozDiDwbfAwETw0dLT+DS1siJJATC/ONVE+g
7Ar0mOjx9kwIwAnxl9oxjvacavMnBKU+Dvx1rK1QGqFc4S8ESEqnm8SRx8SPfqxY5+VU72g2MYZr
pNGuNGf9egPW5xwzhIO7oXCZE4jpZWz3pGXJahGjxe6IEByHwXB80hmFyEo/Ba6X4eQevoGtieds
52G5o3YbE6xZnoHu/hFWinqdB+kAALmMdPUcSv79j0tS+gkWN6qean4iORJdTgWQEEM8gbS8Imck
dyXjUUWppu+gok3FK7NYiVX96kDw9SKcbacCCNUzoJ3cUz99kNkf3hMfJIhZuqwDDe3y2e1rM9Ai
f2v/+/toXYotx25G0kO+Dimrwh/9fbv9mesUcMYjvV6qnWAY662MC0DTt5D6BbKmeYHPCXc9ZxUe
MvLmDw1XbUna+Kq7Yd+8k07R6LK40tbRlXyLywGuzn0R57Z+C6yq9bOb/frT3ipXoaJXF8KU0k+K
HjUyr4FA1vNJ7Svj2wqzoc+rGiIfWNy+crO/Qr9a+YvRnQ7IL597/TIJYms9kT4vqVAVfhwWwUZt
vGdk57JzDUYbM6bkkeGUUe/Fu50IFAVTVq5+Fr1EZgSXUb6lRm3mYE1lSHXqYiwe7PRAxDKu47aM
xkwMsJaKJQh1c5ReC/oYqQpvq5Bu1VCpJsJtQov16zwI/6PEtH4bVzmoPZAVtgdoJdDokZNRAONo
9uFEXROZsjjUQg0qxb/K9VHzVHP7ZycYHMt+Vm7VtI7cjPylAZuoiBhGx8l5wiwfVAk45Fhi0fdw
9fMH6pm6Cbe3XTk7FSAJuFSH1AWr8wGO0Xc3wT/hoSz9Q3FjO77m0dqPKPaqg3zxF6sMynjNWJqR
Qs+D/ccB96BkQdoSLEcDyuadLsgWhSVS+kuUxAZ0wz167cin8Ywbs2qPp/sVaKGNXDTqfhyZa1lc
J3y8cw41mCzVBRUlKfMykgwiWcO+TwfgebtjQRypCgwQ54djVnnMe/ZWwuY6Blygy9ezJnVEYvPC
dpy9uMURDmdISutfChFEfxrG0fPhsQ+Lb+kw6zG044gLJiAPah7pvIr3ZSUTbWZSnhl9W57fnuT4
ganHBK0WBhmbkH5YYZ9BEl/q0adoEKYhutEUmb4tuZlQJwosqLKKgwJQhBlzQLQQHpi9VsAFuShT
RTI8wUwbUCQfWyr5FTNvQXFMyoh3zYu0OhdRcZo0ORFVY8lKmNKgczqGhWCHpUuNpDcVNkIfyuTn
tnMbxP6VzaHPdYJHqeAU0vu/EUt0qBOj7j3csrqzmVG7M1owTo3GP6Bcss+yQ9Ce60/H4zNzgaFI
GldGT4LDnL1XZXoQ3w1dbhqF4AzOiHWyhuDY6v9EK1AsvjMki7TOpMT1w93GGeaLpn1Mh17dV7i6
J/i1+pDWJTKoem22HUtGquCEL3rETVgHMTCA7rEF0miNn/QYw5yB9EA756Pzyw8eIPV/z7HSR9j5
v3zQEl21dMiajDj7k9Rh1kmzRVswCE1EJcQbfl639VEBd9UWDuX3vbpc9lVYtqCu/vCO12spUWXO
1xxMSKW5U7h3V7WJDDcHLxZJ3dXqn/T4MIXru5CkMqglzQ7f0ScHIG5tpQuFONqsc9RQ7PDYy7gV
KkLTWv4DSEyaVh78U2KBRXD6Lg4ImPHEv37FxW5Zbv2iAzS8yUInQr1FT7yPLD8P3JwjWewTdgOm
UWEVbvmEIaMTPZDncnAjFvz0a4nUAS0VmZFmnXwiX7yDPROrNLZMhtqx+luym6YWGW7fj5dA0NC6
dw/j5+Kr5QEBq63HcVY7/U5yL1LyUPpOpfv769yeflz6suSbZ5DMy5dAqyI9zr6kYX0KKHCNPwyK
O1QAmxCie+1o6ShfeAOxCjPwnqqAsk7m8lgq7pTWtN68DC8Q42LA9olDb3iPRfUenFVV0oFHC09a
bXmIa3x3IwfrbhNvlNLdLba/MWZSlnNDGn2soxXTwE6DUeL7zV4X1FiSZ2OeefyBNW2KmPd+gsgd
K4YoQ0aWEmQcWFG7qHoKPv/z+FCY15GYsoaJodCDhZeU5eV/nxl04wP7nqwP64liJ2whLgd8rJ9k
GTJp95ilN/HW3/WcczaCHhjA58gzQJGeXCaesBehVvhpvyH13rDZ9t8wqFK3Wzvy0pHdj7KTSh7f
ELqT149UVVKhSNhOqCdEX2iAYXUcxApmNzeEc6r5P+rEDxrNwQxAEsP/AXJawVEybIL5qxV6iIgL
XQxD9oQGrwGKEAz84Qd+WI473lH6bAucgckg2mZ0PiNQQ2Flnz83x0+4j3EByZA9vn53T+FdP90u
sme/fVVx715dU0z1SUxZqyhPfmOkXklAdMvbVFD66Ey9p9kM1/J7En57zen0831x3QvJXUFg0Zv0
H+teAWqCbj8LhZtcLvKvxZSP2htqcpRsWXFBO5+mfuiplcjhM+7szHPE4O6wB+zWT2o4lvB8HZXd
dtkbWXDjtfjLgwR8TCZT4hho3jaDkU2db3RTsD7Urz1yQjRy7mMH12nwTdN3BYxQeIoTVAxhqlur
VdbYdSaF9My3V22aA/9cRygVTLJTg7YRRkIqGrog1BLFAnosKSyEWRX7fjW5Q6drNWsAmiVFhY6x
Fqudh7ZgF9kaFvE+6JjkXgOjiJ6AleyeGNqbfnpED46ZBl2+5hq23QdTDv8fVfkgfoBCJm4NimDZ
T3APx6mc7AqkTm3V4o9H/Hzx3Bzr3lQupWzLJvNXtnxq+R/XuN7gmrp4P3euwUJJUtKvAx/8dEcT
uHTuTyYbDwifkrEs9zXp/WpOmkFp1UedabDwzNxO6OmQsY/BVQlLPWDYtQMgi1Q1jty9+sKQ9+Xc
wLCZPmaqoJd99Yjq/QGzhgx+mhXzTd/gLvhuMMVqQkizmaADoNid16YpZT9UsDkpKTLveq+1Fkqu
mwNBtG2VfFofFNvoVn/YSTq28ECjPLiVgHmUoHK9vD2mqVsmLQsyZmFSqM84y6Fmt+n636yqo/ms
3oA5rSug5vZi8lWmpyD79jE3DIMKTujuqMIrnYTuZqe1OvPsTcBUtA9v5Mc+EpdD7LTMig4F4ghz
HDHXpXwdv2wWrKbiCLiuykuANuEfYLj164fb8VuNMxb9x1aeIMEhUtBfZ+4OHCvAQsc521HQZukj
dUyqjbQT3QReA8b5TskvAhHtC9aq/wMdhe2tookTlQActtvd88dCMfeBNBPenDi77+rGtMtwgFh/
edHn0BiMingSUiFYsVxSgoz3N/4cypBbOsF64BpTMwm1rzKzF/MtaORMwVkQ/g9ZDKWuv0lNbmLq
TiSzZRK4Qjo2oOyeQQ4NBnMJO5ZCg31p12spNRuCGivE0r69cm9j9DWFz52udcReFnT7gOeqLR8Q
uIYqLhNizwWlic8aoxCfziblQnY4rhT7FjQ9l7gx3MF7oeWPk1o7JPCV3ZTNbz9/iCqvkdjJEqs+
gyUFdQzY1DGIxMGKWqDVVV8ylypOR9QBtOMa7a43vke66c605it2liw6frjfL85AT32jMfQ6p7vG
7S/f46IG8tJru3JWMePtaErRI0NqEVGUn1Ykh+VrE4pRK5p1IuRabCzjSlty0dn8+Ywaa055nQ8t
Eull2LJJtt13RMT8zu6y7lgA36XkPzz26WHmGB2KwZNXARSGMsXYj70yr8nBij5d4G7+Ahf6Xqre
qE2vVmsJrl6KU2RGxSMZHKHiy9ypBk4rHX3uNswuEjxPru+3AZmimwk5copkar6u1kG/UMf7YcTc
AM4yC4PGT0TGjHcukVd5UirvvKqhum50CmS7aMdHkLnmgegUe/BQsEYqujHc2gH+Z/jsCKm6x4My
0TUL3Unvor2ZFzVmyBn0rxbGqej2FVTfvsqBqwwYp25WCcUoD2sErjM2YKFhYQ+LnlryFlzwayv9
XbtQ9Wh9haK80e0xyjMU3p2RCv9yJnZtt26ShmWj/nA4PhhrhL+LPa4vkODvCWgoJlbix7fqrYoP
eFkcLmf+vgPKuPE2t5Yhnn/iqdccJe9Hm04DvD9aeQ/7EACfqleAzrpK4xoTz3PxuCUlegvPHHWr
wuJJekW7x3ar91GqTUktvr3aSEgv7SaiWuM41h4NZuZ4+6apQQ7QVXkxYMClSk9mscoWx/IF47oy
KUCBmMmy/4d2hFc19Hwaa3wtFLFSX94kx+84HAEnJZrwnrWFB+jhCND2gZN7ZKvICkxwikQrXlKi
3x1MmthDKclHUpqT3sk2GgLQjj26ZHPQ1ZKujmcw3I/8FeGjJwXKDYWrVhOyOuXujPhw3ca46eQP
HAlLFYunxmbs5fNr9dq+ouNudNTVlPDbrgzdKPq+zSSO7TxUKC3oqJCK69n+a/OJlTD0wpTCb8no
8pR/KRmIGViyis17rad68tMwI+ZROx07w4+dROqTJSYN5jKRWpjTC8yZrUDoOHRpYLCpfBCJX2qm
bj5pIK1Akn3DGsNhSPmctKMSaX9NUfw1CSrn7C0xLsPxtfqcetw1AmfdXc1ph5fgedYvPWgpYRcp
8yvaB2rEIpGu4/ulm3fT6+B805is5m/9dPZ+jfaj7WBqQgoCi6X3xWqJfAJYmynt5W2OMcRCyk8u
bv6UvoV4IQ9t1dXUkaPb+AsO0nwxw+3ASRCYEsGFkghrJFZUd4RaihIBWlOzaJs8trwNEK8dOZ9v
K2BJCtzDghF0rOI84t3tKIg9+DpjoxpRGX8oYXhSsR8nJjjTgSyL++ssk2zT5n8od/8+OxPElvS0
p/u0Ifw3L0Jl8+vPv0LG+voxBNICv2RDyckQuiwxdwQswNf91FlVYW0FwtJZFXj/nFtxFYm+N92p
TUU/6wUT/ymecGI3gIBGAM/tTdXby57X4HQbdA9RwrZSwberpL8rqnI1LjJv+wxo+1yZZlMyVy6W
oVfYdH5iTgDeZ74GVfEf35DhDTupSH5iXev0M4N0xcCr9zgHnkm9Zo2h0WX73t9gh4EcRVCk4sci
IcU2hCULmoSURXYsZnT0M63Ajx4g2/aNY9f1app6kpzhIKcnYNvA4VYGYBZC94dOLzCsmrcr5xFH
9Q6MtwjzCuw4avcFK/YTQihG5HmAlUjTwqBkUBLqFgKIuetY6nwX+OEUepfA2AlOc9KaLB3NukXa
Ag4prFoGAZtElWGA1WgrzN6Scp7fIlrWLX1M8KHg4xLPFo+P+cfPSpPVyu7PIjJItOZoZgQfyHr6
pW+fX4Hv7FX3YHff2hWzm+GmUnUTc3xvlCskMbPJcDjTT78NShS843PEjgZA5H+3WEobz5gxNUvh
ZQ6dbD0gkXPqt8rknWlYeFCo1WrEL70VCViUHGsHP7zbt7hh39E0ut2GeD3GyZ/wHeZu/ZgoSffK
hsjFB45m18VQ3IjlCjxR6X5yRw23EGZgmpxbVxwL8NyZuIlUdoOnT7CeWTh3R5eT32oNfrfBDTR/
OO+JxA45xgUS8i0CpzJ0xj1EgCLPe/0fdUPrhCOB4QOZSjh2mWySO7urIuyOPBFMhHTW7cnTi/TL
8wMcrtlST61RCVL0BqXku/X8KKkVubxl9T1he/17gHWjm7BayqICa5tNdD/mTIzYGeu/7I6lQfj8
66NoYAA5J/fxS6OHgYJn/YErjepdPUbMFtCCvsU24COCw5VWbIEcfOsmx/UUQgDaU1oAwIZ7IUqa
XP7YqnuUNeXbbOta/PyU2mgMdaS0mT5VYBzlMgtluxSDsJkgl1Jt0tnh6MQuaYoizSv5UbiMfdVQ
mAZsjnNNlrC38fFgOl1PD3HV4Ysymy81KTIZWNEWb2jqnbH2mKof/ci6W9nTWY0sFIvsYMTSEcux
rW/hboYvzepuEsero8aEXUdFeUP98cx4Ao1kRtrYc2VrsdYy0i2mgLBTAtQECDTkdDuYRquPy4AG
UxxmYxFEUoGcfc8jJQdSUYQYygC081r87nn4q6p8qV4n1JIomhncy+lOnOKdtat0LasOGlJa0seO
4yRXYQzRZ1pVUJ7JQU06thlKKvu84RlctxaPw3kz0QZOYpaQ493vVxTjH1zywtyv240y3rnlHBVO
MUU78kD7OQgZfk2UOONJ8JhskPbfJT83WZwivEFCJo29xQkJLH7SH1n0ZAPGT3HbTLEU2dIMCWXI
X+w1XZFv4LQ/WdI9iyNroRTsDB4JeNo8dJQmQF1iH4oZ/92+z4Svy5fPpS2ujLVKFfrfFtdUy4HT
cXkTBEh5pQrGSDMuHKAFFw5MyN0uhQQoSbNxB3VY7vJx4NNgVZKh607W2+IPqbYQHd7qmm4/jGdo
oMgGy3h4smV2PHDOVIhDx1lFnxK2kRShiSD1wSI67qNM9wPNXc7t5o5UJN5VkcnUl7RNn1AHRJrq
XqqBGEQC2L3zBo76LV3wS+6LRI1R1Vr5pdkEOx8OByxrPSehse5vucY7j9QRAdwm8F1r4gvqTMyP
iBV1OCHWcena2vFMJ31TYFx01oXVCykZQX17aiRsX2CQLQkp37nAoMehjRytcXvWMyT0sM55zpmp
PoGL4ZKx02nQXwO8jnR+fLROBTd8z2YH2+iszsDTVTn3xFeSOKrQY82h5dAqjyZ3szYVRYolQaJj
bvw0JSBG8jsDkwc7/kl6OQ0cQ1sM+xQSKSZqCwtK7ND31lOjOaBbYVMlW2cJP4mzFchPpj4ZpjQ1
X5LU8SMCKhDo4A6fg+FzJFCsxJ3DYlfpvy7H/3JCv/KE/n87cFLhx6MDufPvx1sFb8svicAmRCdB
6IeM6ayczISq0FgnMByCFmlc8Z5KG1+o45/e2kfQDs1c+Ol8S1n/KSuR4X9ETANZMZT3+P8IWWcC
/8J4kRv4MctAUW9fEwyQ0pB4bgwVc6IPnK2ngGVBV4InTr/3Rzz+UBO2TIjh+9DLmTXbTlFVqcev
W1P1WYxrYCclRQTo6OhjbgWv3wEOgfTS/7/ZVw3ne0F+MwbQPyvBT2a6DApqf/szsK1yZjmQd95m
ARhZHsJXj3QF+VwalPG6FYOkxJLsHIGVO0D9CzLyzCJ4bFPLp1K8zxUsFBKivg/ZpLf0Zc//mgUw
4uJY1MXIl3Aj5qA7FYZgUjtB4qstfruDmm01UrGCy01z0Xhu/7KPQUF4AQI5ZsSb+j2UxEoCQHYH
4xVH3LNxgg4X1vZCQeUxoq8A/vDqHDAelK17gl5MrgsxEWSLEMetXeRmtiNdiK/3TTk+1gWFKvCn
brZQrWFp04G0M+fs5agC1O8VXkFFquXXKtJZudOr9+l0dSB/mQAqoGf2+H7H65auMbZKXxWHXX4j
2dh6ZKxCJcQrTmXRfC78cm1O3qFzTD5lEOXOV6puiTMC6k8nqBrDl5171SCUNC2xDskM2ZFta6h1
Uqw91ZkcwkYJKpV0UpLa1dJSyK2HsMb3U7eXW7OA193oDL+FFHJtmlypF71ALFrfuzH9LK5atS1Q
qquQ/ccBm2CbNRFukvx1oBjoB1UqaXsHZtQCGf8iFx9AlDeBJonnWR3EqvdPwDg9sp4CAI2RRoMD
EkYK6ILUp7BSlCk5mH/3XyRbwMTGI3d1kWnqmI9OFHY8ZrOt+uqcEOzsbef2gBQ5tgXIVL0oFatq
bDB9JFIV7AnZVLVEWX5nzmf8pZ0QW+7HJvCEhdKfAKt1JoG+xYjsLTeIU1osS/gMLYfGm/snTGRY
/bccYpoVP6xuGUFkf7SGNybRJ7YD+le5yK8z+1YItAtEiARmqPN8oXXZACRELfX6nb/rqXxKf8iM
D5XNpR8ox4LPDSZAfipkAhQ/C4Eow0d8f9ZhU3gSJQ6YiVj+wxVHg8mzcB5CsWIpL13i+ec0Vs5Y
pMoxlePyE5F2tTpN9VhUsvcfgUJS7zfS5m2L4c24iGtZDUvwXKFon340eI43ZkdXnAfOmgjmePTL
RISC18H2GFZT84F5nwqxqkgL6dYxbdGZNygUu9aJSQ1EsYQ/52ojZAXwlSYPat74ilbWRt80MNtD
OZl9VHPvQwUNwYAMVLNSY3JK3ZBnxdGjtSSHMc82tWWQXnqqD0uxqnTdJj+7/leTsIJza47s8JV8
btUe+RrkhvM9s3i8FJ4wN5/v4QSA/oCC0A0dKI9JxFJlDdxbtO5jqCbqOra57ItQhuFA0rJNHihI
Fg66GxoxROfUK6uh2v5kQoVRicLj0ioeDcFxBDp6TfYQLQ9i68YLKXhqnZb0OZijqLa4AEOoRnil
rCvqT708kE8mtqYopJznpogfHpvbaUg0DeFAGjbJmET+ND1iKUFuUPIWQlYVOj+6rrh50doL6/lO
u5fhdjxmEImlYOTqad+11jhkSqwyX5eLTU7CLhMOBESOlS3hZ5saKl88yYFwyUw7Ri81S+n74B6J
h1H825UFm03EGTompGATC5Q4BUIC8kgRr+3x0whBDLIppD2JTp1ERhUtfFQAWGeWvH11wLfXKTb+
XO+SPn5agIraqD7ReT2LfLBQF1w4s6W9pBVqIGGAJ2S/JpE1Uv+xzB0k0jbZGMQboGeoPfaXl0HF
gTn8GOVCZIizpUu+WzieG5RJrQCgNGRkK1j/VDOI8lYC8+Ym4xXfEo3ODa5Sr8EXxH00Fp2BbgWo
pxA0867PSpU3hHf7TiPElF0uSvDe4YFdmIFk9vcO+ok40j2rUXhrUXSbVjTDIYHB+5i9KiCI8Mys
52YlGY09HE1OrGM+ZTMra7m0vjdmKUbkPdpnEEE7llfU8sgEwFDvBR1ESzLVBsAHTDqncX5QQypp
3Xveg38PvwBb/a5Wh6+Eywl91CmpAf2PANEdfRe4PP9qTnc5N+Q5n2XUKE+H+N3dAl66uC3TT32s
RpI1o1A7X0gGj3EsrmFSbuPAR5SiUH5ZMuOU+02GE0EdSVP38wt1r0e9U84UB15CoRXhUJi+vi2w
JaCm/ndnC6EN4GG8SbyPMY64TF9GEsoxHe2LLLwGOuDb7jjyPUhzsBBuhcIM4ajFOpwk4kQqQETv
+e2L7ujreoGJeKG5rD+SEXo+R0G7BwdZbJr2blafL6R9sQPz0RQAHB2DMieMbiFQOvJmU6AMyinC
/XMVOIfJ8A+eIx55ODGlq89XkOXrBGqjAeT18eOrQiELzUZ5G1oYj3RpASML95W51INxfilyxibx
qVVs1TW/QbeJ9y0OX0+kocLLOyaJLqwzPQLMPahDA2aNlaxLPpG1YlMsiqJ7h1tDJlHGBoBaaXF7
1G7ic5Up3MwztBZaH5Ch3SustbIcVqAfzXQdiE+3QXIDhPLHH8sOlI78WQS/QoSw8duqBbvRSDQ9
WLwtXHgSrYqTcMUbpRnmQxJ0f3PIMo91qIMFpB8ojdWW+Qiqg/UN4pDBO7yY69p0Y+UsBJewxim5
7oaMH9mXFXqBfW7sOvBEsBOevPVdWObAwis9w1x1deOw8wvtL8BUEJ+hSOmrezSp04JWfmZc3Cob
5e3jkIMEdf9cMqYXsz+dWcJ4dVeLaao0kSW1R+ifgo+XHryfpeTevKQUDITfvD9NXKaLuMKN1TXx
cytnRgmun6sn60jSLr5h/HAiwnMxKm25YHJYbPFYy6x54GGgWH1szhmOypNgCcjTe5MufmNqG973
ZewTZ0GP51h8HiDft2GffnlSvRIyGs8mTFUmVXUCuJk3l0no+xIGRxejSELDI0yVtNFYs5ezzcST
hDsJqDkbgl9Zu+Wnvb4/3zkTCJiYSjCArSKRlYBMSsQr71/JyX7jPx3JQCoQtM+ze9XdsiZhccJd
i5JY+iZdJPt+ded862YDb53V3wTLXAtBQiCDCh4h1OgqSbM+d4ZQ1kqE+NseuLPFJYpzLTv+gV2Z
oJEorsdv0Zd1CKraZUSBFZ3bbWwbmzOKKvoQngaNT5ZktOw1Q4Q+a6uFkciPf+rBvFOwIjKrlFov
IpsTOQVxwWYv5yGpIxSsshi//yevJ94OQyfpyf6pgQwvPowP/aub1INI1MBYL17w3oYwbCqYa4Sb
CtxfTejVEC4CcwgzipKbOOyzifNzH9Bcx4uowpQ3ajzhwoJ0dKJVAPhwMSMNv0kxwu9jrROkock3
dRX4v1t1ZDZ9sf+bydpZYSugUd10wrQDhD6F30eU0by4q3zUKD6aavmEvPjyyG5MzJiFB9/FFcJS
+5Gc2bG2OAL9FJSAtXZxF5HZOpQISjdJvjYnLw5EWXj+D1bZUwkInZCduzpUb2ia5pTgnPuG8fHp
vpgzrCuVKOJx/FPvp1AX5JQUoUxcRke1TwH8kD/m/7r1nf4ICdE2D9d06CS5mD+xdgCNZf+9OGQx
ygSTXwDFa8gByoNiylQHtFVkJt0x7lFm4mInJo/1ZJoyNvT3+AUqnIN/IK9j/BUYXJjqK54thEW+
mck+kNNRW7bRbWEpMjFOl7uImjfxhymqefTpg3fAHcPmeNGjTvSjzgB0gG4ubUW8tAMTNTVSlKqX
/ZuJL/1OzonaW6mPqGZQfmcb6oXeVGkL16gCsU3JQHMu2zNp59Z7evpxqsekvsawXCKDigUymFAK
8yi08yaooR8uJuYXvRAK0SB1mvdL1Bw4nKZr/2u15Efgosjw/Kp2lhwf3Rv2UVLoBd3+OPNJX+bQ
6ns5XdmhXgLJmcpAw2vzEpC1/rZnSRxDnSrxeSpf/rcus7VRm/JboXYxM1jsg0JFE7lmf12tXtl7
m1knV5+xXHxeiODH6V5+M9iEHnFVM7lRdYlSkFPtUpS1dqcpk3zPlnwy+HG5/62M7EsisrG8kspE
Psg+jw/ql7swhhVQVFsFCr1aL5tCu/OlRuSkuK1k+6OaDGUYD2p/fbBbnsgV2eHTKgMWsh7vadrx
zp4W3ufDwBi21sIHpw5fikJNrYqgl3CZkr/YU66CBcfhv3tsWNoKoHO6sjuTn9w7igyTNzKpjkVA
OPpku6ykP36yGaiDofBesMGyLx48pp+nRt4WV+Gyw40Pfs19h1rQXSMC1CdNk/Xv9sUkcODwCery
Ep/r3NfiqW0XRYphlQlTrdzAx6pB1WNiZ+OA52MJdLaXUkvjGrpHLjpQmoL68tmwZ2GWqUCa2l2C
7MLg0yNRsOXAqMWawWHAgHGbGoPxdwQ7tOIGDPQqJHe0T5W2UHZ2Uy2HwpA0EAlp9KyYBw4ZtaiL
/UXNQaEuqjfSjsCk8bDLOJOimFd5qHC0kVEs9DqEfVyeg040DBKrR+L69nuLjcDUz5SgdW3MMmNW
x+0Q8CPTIqMygK0Qke3R4vv8ycsLDkuM8g8gdPZm9XgsKLoEFoQCEje3/SZPDL0CxH2aaLSAnQXO
cwl0CBRxmkcwfj2iLaSYtWawhovBrcp4NS+hvPyht+awtgTdasRX314RJoUnb13UKUSavS/62/p/
CeyAlc1NM38UuUN/Ef4ld3+xKV0W7uuwg/8cvTzFHKQRYso59lNMKPS+dKZ1n7O62SZZzC77vCXm
5WJmjXqJgWDgGzEjaKemQtm80bU054R2DDzPliWuG/cugIPo6YhehXv0ugntTYwn/4GppSWeoyR4
JxxoZZs8PKCn3O6yiiyPTVJYZ8X7MAqdCV5uZFm4M2eTUk5YNaqeOXjsvwapIB1qynrCgmdVucjZ
WZs6NMFgce6CanK18CQqxX8QI545wLhejx5NiFlYqfPKRlVWiVu9ZgfbUbRpvFa40GDSHtS1J1pZ
jkHeUC59ZtyU9yDkeKZyXG014pcZM4cA2nU4Qxe7I8l7gUU5i7ha5g6xZbb8zFV5+tRivhPyVi0a
Pfafh2op+18T8xLOz+unqvpRi+6Yymz1uda+s1/XmolJ5UssExYFm5fEQ1VqebrxYh8M+wEPBNQA
tGVmvzg8dr2QsFAPJgDJmrV1RL/t1BApyXJIGZO+9sssDNoYtwmACANuDVWpQyV1a5aXXOzgnyu6
cD+heopDwfhXtJ3TcLGVB3ixLTZHEOt3XLvm+zUwuXEUOD2yXdUFooT5KikLBU1Kpyi2nzxBHRTw
0rmLMHuL+4vi7c27L4w7pXWlhjaKK1hOYTPopbpoE/S32/9u7pIYlcirUgUUo5xqJ0e7f4lCUJ7K
MyqdpjiwDGoSozkJnnWvcXKJ8pNeFwU9lNjG/lXdmxepB7IbgB1BOBvGSFwBjHt7G0wO2wwmbfbN
PGC1F1IEwofkcrTTlQ82R537y4Lr2IN7jozw93ktTqnXPAGFa6Oigf8WowvnOa+BorRCjptwKxgX
09KEA8w5wD+CHICVUxsio/Ptzvl/6gz7nuWBkKAgrlFesf/gPKPB8tHt27ZPhZO9mUlosh6klz3h
3W+zI5Mtzp/OyYqyvpEx5Kjo2A7frBD8M/Q/dt4lmAig1qsxU37ug8eMz3UyoBQIcMRnPyzViLzR
9zRVy+jkC3pn9MYrKEHmfRNJ8ohssyX+dlN8tQevEe5ydw+FwJ7C4yCkL1ToYJDhLN0MdeT8yBiN
WeV5FLo2ibuHePNCuaDnYiEwt9/sXTESvmf89tU4anQPR2We/wloFNqE1sOlwzyYH7x8ecyqsrOh
m1X6I0kc9mCqvbNIWgSrsVLEF6xauO3iQASJRYL7qpzzfhCMjMfYZynvejwDmqeoBOANmBhy4aXd
gTTReC1f7N12iYinGElqgM9Euaajx9QXtIfgMBSwF02kAQCI8US8KsSCAwmaXIXBnt3rmwRdceTA
Eugla707bLLzRTEobQb9e1bl9hXfmZKm7AezRXUkp6qhJDpvmKNGXXjoij5q/+5NE18Nc0yev/7c
beVcIvhyaB2N16xXGKeTjYgY28jzCzQch42ZccYpZdvBJxi2AGdsDnEP2K4ZUlAgwZvKi4B+jOdH
yP8IivNoS8p+XGXfwhre7Xuh3vXXD8lAAht3BM5C1nKnXyN1o01iCWME6FhHv4xpC5ErPrQ0a+cA
+0M8yinxCI+Uwdw+exzWuj6Ca4zOgRUCxzindu20z6C+3R9RlYrgfBnwxoupVdvqtT+sNDNxNUaZ
nb9JP560zpuzbwJYJs/0acEeB+lNe/h4h72H4TBSqWpsQwnxUb92S0Pb5n+miKa+pv/UCgsnKDFu
lXLrY1mXo9kVotHvqCvaUZCs8OjykNlRAJAU9ltDJqh6m55Hz7Rv3dOHWvCnYnrDlRZDN0hcpAST
4xDZxuVm5lNrEdiTlTHqQzra37XC9GuyMBFVXprBsBha51tjRe7O2nGZNprBcL5ulN1ve+JASpuz
8SzLX+pyqgkPY4gtCUELntNOivXhAbqzsjdiSI98zrGyD3vYEaiVWcgUD5pUn8JzwcHUYIUQK9R7
vVODqOpg9uLM6oRDx15z1a7mkLQftgyaICquZstAPaNhTzF6IRr7FJJlpnumM56MgJul3RZU1Qe1
37smb5b4OPwQfWgXFy22F1ZGuvs1PFX+wwkMpw+hFgKaUs9KWxx7q2t9tCota6PhrehD+whm/+R3
ZUbJWVijxSgmckOseWIJVRBzwQ0EPEbiR+Pj0VhGoDIABxzgZSZyUvbqN8keKk5WKtpDui+hdykK
8kyrZ1587Odj0cSV0yeqDeKNGiP54CU0nA4Uza7dvb5Vx/1kFW8tM4tNcYk+LZbw+kXeXLOMz8bz
XUFPSkTxQ97jnBJSlp4azCS1J2G2TpPkDrlzLALPzZWYuHbyrSykqiMEXNIOw8pzpkXNFlg60OMX
QVv9x9G2QyQxzIhvV18/NcqdnzyFJhuAMmY8ULAdB9q/o0gBZfjymyaz0eWqXVnVodnK7XQ1QeHh
0nujo81KmQbiQU9TytawwaufzUOa7FZnRjncwiwLd88mFz6yk66SlQio8gJwI7S+xSP16xOkRkqm
xuUYd82LKXhoXZ0wrrcOSSYXETavBo1C+NERW9WT24/mdSXN2vut41ZtDx8okx/WWD/J5FS9IPvw
mHVhZaAOz/nT0SeVddhb1wdEdKZdDxFROTlC7u8HY+RC0iscWcbyl8T4TRxcRaSadT7AluOkviO2
Lx6/mHil6jcfc8ivQMzXGOE47P9CSqaJrzqqU29K/F6nqyrQtRrVAPilF53ZlpY2sRx+nr1lxVoB
pQKgnX99gmeZu8m2Oan0EWAHZ8hjRGqPCXkrtKWmsPfXT1YVcOT91UGBqqvgAL0ZR6U58bv0f5e+
q/3FU6spBieZj50ei4Skcyi6iUHe6r6WYc6dBO8OeOAbOuywNTOChcRnWfhJv8l8yrQMZryR+h2n
6EHet1pKDVM8ObvN3PVhUyGf0qt3rgU22/PCFya1vi6seL7YlU0KUxm5EoRdMPzeCDEc8x79O7JR
P4Yge7U/jKnNt4p0wXbskQcHaCAdSP3ujFfubRsx9sMkdnT6UPnES8hNFpJBlDOfWV4ekKb9G2WJ
qu/Qt7A++LFp9hoG3dOAZ1JQ+3y2apA8sy8i+dnL/FzzFjY0NoTK6ss9XojOrH8MOYlZIRC2rJMk
SsE8nTDQax4TbwvTe2CTNMnwBquFI7XhCL0+Kh10h1tPONjYtYPI5fvOoPxZgCzOo9O50lReUK8g
hRoUaVIzznQQUIaQa7/8sZbvXciMERhS6QSN4KFAZMjUdcBN5hQAai8YIGoMtzrZu6NOHW0203HG
iw1f5EhGTEJ948KNldRha1wowW6octV35Rad5gXEseZp3CdLSvFFB/kob3qqyGyWYGwGn0zBfTFN
6JDKPLaeDCgJD53unlvnS6bJGCx9dGqEKgBRy2sSOIvqPmdHRrG6zLEcuen+0NCDTuq9+AXvJnFa
1CgqrLHp3LejUy/79trjLCiIw1bVfV0grkR0JuDdOSR/ZB8d+mwtdV20KuqThSPhTf9VOJzDgZxV
jE6mffKB3E8esd5lsRxxSM2bhR2L0lIVzPXmpgf6/V39CMRWARl0Ex5B2uLOXqAbACbuwPbxmTzt
9t6QW8UbKlkN3c7e7JyYZRtgtygp6cZB3uJBjhgDFLMmtjJyufH2PfB3+LnfmIprR/xFJ3aRJjqb
zkRw9wt350Nnp//O6PqYwVw4ifdEniWt6PgHY4gqAvRHdf5S7unNJsy70uVEIglxLti+/bN4wBFB
wLJbI1D2K6WDMVHRHLA0oMvckKQ3v1H9faL2yHym9MIHg+YeIxgqvk97DEuOS1qJw+KLgXMmw8T7
osTKxsBEd+zx6uXhDJLVzQwepNihnE5niOYodakAnC8fJaSU+5UgnejwR67JFqWGn5SYSzwIVRYV
5jOZI7NuR/RPcYPOknCHU2PJdUKqL3meldlWAA8ydewM0qwlWpjB/7fw+alqzJCRPIJLMDYPHECi
yXemIhnlgIbHj3bc5DUvfri0woUkXVThWtXezi3Db3NMgDXJDnPACVad+6YLA5Jtx8q3rm0pxM84
PQsMfJTAa1V5p9hIzgdl7bHkDU8X9Ma0pUfCFdMOKkmWqO29Gi7tpuClwKXpLlmh1kW5exoQF53c
8BEDUDBuI+VqbSgzRPFkcvqv9GiEGtp9pzVlElf5FWIiLyG6HsLvZ+mz7Sm1chUxt/r+4ZMg4snc
oXnAUippIfl4ZJ96vy0yZHXe37rLap7jrilHsv8n/WYUtiVEAziwQpwo6QQzFkPTcVgLMm6uUiz1
p4zFizIEF2yHstQtGpBxJ7IzQTQJqyZRnpv9L8OlC3lts3L+RSfun/liRC75i3aapFTcnlhHJWd5
f65y4dB93R0+adzvRc+SLsCProhD8BvlOxAbGnyd4psUANyQx/9i0uzK2T5xMENt7PQ1pV+mGdM3
XNaaMPz1Q8cEO6cfBymy4Dp5bd+C8x27mPEkdWQsRhmS8ehgyEiEUqsj/OE1eX9KnzFTINR0sm69
HuAIVadibJHhgmngMI69zIv75DhOJTB3pqtOl94PE2fKMKkXNKH+Qsu/qrLHrlJzOiBvzo0gcv3l
OFg5VxFY5ZZaDkuRC8ekw2z+xsln+GKrAIsAeKxFMJmtY/EwXETURlYROLi9ruQkZSOpimjojeQf
GoJE15MupBcF5NabpTN2uTyh9Q5PGo3eQJEueh5s390i7QHO8UB7h2e42c6H+xOziypF9trA3wo2
IjcWcIkphLSUvPOyFJuquIU3tv7qkTY5OrJp53xn1xh9W0LpxMwDSlP2zFT+TH/HTp8YfQvFOeQ9
LXUHqINUqz4iZ4nQ1QwAwrfsm0ckoJlRBVDg7cdNJYi+/GPEZeDmIqSPAmvnPLvVDFq+Vrii4EHB
j6KdEE1sV1trzngtEYk1Ezj0MHeRzj6k+Bvrf4YKF32GWvV7IViSXR0GP0l6hmWxUABLvYTExLK8
e38O65n01F+xVnVSCuL6W7bBue+YDPRFcpVU5wt8k3UtMpLMaG2Icgkf/cuuR902v1OVyzyGWkNS
QJsCZ1Dxz+IFeIXQDxbNLQOReWulnOW3Ie3oQy+UOOsdPkpBRvIU6ufYU+eY2geJUmnw2mUoR2+v
TCKxaYrgJmwgOFbp3JaOG1j5LJk+lL7tW53ufWOJEVsBmXl7lW7GYmIyMbvx6Ab0+wEHo+/99z+T
rELoo2BYTXLoetiNS8pNlmGqHhIMXeYOZy1ICGaA9y7ZZD27IV9TBHMyU/cPoQ+OgMULKsdrQQya
L/P1p74ej6XYPNIkv5nXIJLuW5skhkBP4AOmpexcSwrjgABg0pZZ3+Ke1iu/3uGieN4X1Nqk90/j
SDE2FAb2e8QvHuEXqTq6UK1mgi/5Nflo3taxs4gxj5Kuze8QwYVHQDfy9Z6U9S54JwCKiEmDDfgT
3Is+7nXLQq25PUZa9MtozeK4xWcK+OJbHQhLpjtE8xWbzj9ivbP+qxgEUsAU3DEYxLxT3VDiMd9n
2VhQhQj13uo3635Cy1/262Wby68R+dIQyAKrgr171ajG5SfYn15CvSrfgii/fqnwAy/AveIrarcc
4GP1Avyv/wnCx+h413HMzt2+5EFLpkRPQPV9iHS8T0VFF31VRUV1Dp+cpGj05M15zav04ZHWLIJ9
PKYDBaZWTAbotqN8Wow/mtbiGuoHkCNyDgZUqOw7FhDKZ9q6n39Rbtnxu0Q1QKKgX6mmC9FIrndV
O9igRKYDqWY4kq9u8jmofBmlUXL2LGU1OKte5pix32/wln4I2NVjDfF/9uJjfeiFyBCll2OXXmKc
tT0D2CSrzPv6D4x2THf6pNoGw6nGICeK6+VxfbbJzxEJ6VskRd8yeLwkYZLr0Ul0/4YoyBvRVQID
Q4UYu/1e25ul1y0LAwx35jf9yyBKsl8/z77fVa9SeYTeLvN6NirO+6HdJ5RKlnrjUxOoOijp4YCa
pyiXR7B5n+ofC01GdvauJGzWdj0ickhFdJIFf7JsZz9Qe2SOsR+A0RVEUMRPBRfWPSg4iPIZ1vOj
gnjxKlXgXkKQLzmsOq8N5W+s0DHHU0d6RKWoy+JJZADmdvpKhpcRIC5gmfnExtfMgViK1UKrExzD
imBNLzMWE20qWNltz3G7ndya4y40x5x3+FVRBYXx9mcs3TGi+Fr+FfUJfWEimBgayzXJhTYiJ0ZL
8qYASxihaWimPHIZ92Be1llwldTLB6pZXbRlxk8cKLiGD2WmD+n5fNyOYv1sXlZVmODT42f2tORr
B6Y9QKYIzFqctOGJrmxajTQqoK4MllZnDkOPO92VvR7eWv/ZlcsrVIg3jBxK6z/qBw1PMndOz8XD
XBW9EA5+vc/OosHHZCbQWZhTHSilOIebta0sWKr3QRmFdLuZhhxqVG3+jGcvxa2LgUXwrPKUjJa7
8WA5InZvr54dEB6FL979QUPVPVxP9Ht6kObtm7rgbJbeZV39CvdihGDTyQ2iKGpLaVt6og8MIFzU
kovNvKkkoi88spfRQqnwaWO8vihRoPqVMG9/MmT6D5YoSap09rkBJS7jX+AE3DT1en528mLeXnLJ
uTR9JGda07dQcYIgOkv35VCLxA/xEYX4llHvMDJ6sXJpR6sAX6ToS2hr4Q/qSIaXuFYWJjBY4Nem
vW2s3smMrNpOWAO5SYffN7PvOlXRNQnJNaSvh5IfyTC1KrqMcloy8IbjqCBOYC6a4sxGuprtQrxi
u2ZExZyHOU1IU/qFVXA2prc/FhyQ4frYlC3OWq27YP1Zi9OFTzkgTqnw28pxUa8g5wwkWCBjba1k
R25SOUdOBKaClNeIKlEvu8CkzR93KaAoGDqAB2RaNx28u+BzN6jSEqPRqWw4/Q+tJ2AJe2qfkfSZ
AaWL0yhrGT/yaK6sEav9t8t6BQ+Br4KqQuSn2ZGFMfrmxsvOh6tpDxN8ovk8+6ms/UXyO/eYzjcw
yt4v2Chug/flkBUKjoOI1wZ/58tWgP0Qli6hnG14ZSlKNWPTl9nHUfBZUoLSXaidZLQ6Yj6epwJS
wsFBC61G75TCDY7MM+uC4pZ1ANMO7HmWJoBHlaD2Y968hpnlVSz9ev1VlN234ht3d4QdCbKLDYAF
vfWTJxM5icGGXUjkBThz9jz3RAdW4LdmAEU5c3XnsZzBi8YkI1W4K+xyWdqWodgbmYn1QVuXkMBh
uzTbf2pUwX5GgoTs9Ve8p45eHsqObimDVCwpXwHDGMtTDOIIeZ+CTUbEXqXp55tPMBl6Zt1oDlTy
r5y2V8bRwRO0u5sMNkogs0+RcqoBO3a2BFbH7meHtLAjsywsbisAKwgQy8iOEMLZmVkk5T0AOgh6
OXBL9wHWC1/2RsYIDOESE/7HdmoYuW6Ct6eLfjgmyoC3RJYCvvc0HJArQKD7kF17afLLp5LVUOKb
sbygclt2RcO8vwBoAcrv1Y5y/bQ2TH3eoDyjbTs2BkRVgugKhfqnvlPRTPxmI+GYrWRpjtv0KUK2
UV9eVm2i2+4iUfgKBPCvM7Qwi0iLRqEDyxW82S9/UtzcMb9/QXMBzEbwKVxWzo6B0wBb6BRRVleR
16jtv16u8YttCGiyCvmVnRmVA83Ku3K1cJ/WvkEpeZQgyGjtcSkSmHRVGgvmqK9eSeDOEqhPwdRR
QYVGb/MAaZnxv7F22SeVCSVt+4lyXTGj9W/iSadMaFtg7rATw/Q8FuyeUeHpm0QRN++xBs4ubFl7
e7y0yqHoSR99KxV/h4LmAFr+uYlG3ihsjDDd5d3e/qg0xkPZJP8XJz9EgAS1oy++8zPeddGBQUmX
Nptp66NliuT4wrtUgXuGRtaIyVh7TvExaBGB5Ynws6smWLZbO46uQb/hsGb/5trMQFcjN73HUMz3
NewBPbf2Nf23bmLCubNZjX4myhEg24sHV7FfXulfVmiaMR5yqP5w/rl8MMtWsEwH96PZDvo504jt
2E0tu0x0ojVgfVEXcs0a8iYamho6+JxFzmv2MPaXDQca5Imy4mnwE/MXok0dABqwKlu91VRBnrAN
nJ6Qnp8rz0f0ZbiIR+NKpJThgXWvuoRtckEKQNfzpsAWNuP9pGoYlR6dcg2wP0G92GyOlNnWcp4X
kxO5Nxck9h4SD1UF+OCoROfIBd5+3vtmaLooSM3nPDU4RIPrcNRFrSpBXXVkycV/mwaNMRmmKsSs
i6N/p7utGT7X8ywzCTP1YIxq2HclAq/bNlmtZlVFDzump9XVEuGd2q69vyMXljC3sNOYFssPda22
47n8o+28td5w2AOciP6Oei9LoXyAA2InKWZv7u9jqoYmRqRaxvVRp40VHU6MYY2ZYLgdj78mqjo6
u491JuyIFgLbYqrwR/J7fYdcniw2IJW9urVRmRFGXwkWZaTIruYbU1BKfc+0pINnWZyEFg3h7eQ6
kSmG28RAVQ+7E+SvomKdFRoEoJ6n4G/69AEOTYbhbunCCsB+nZ+VYdKRe7zbujMkU4WhT6RiDmzP
F1rdXID30gzc2TbPHuIkv1m0ViV1Fbcr/GXRPd/ODC+yz9apTfUx0OgbMSgc5NqKihILPszLFZsh
fHg5ox3OdEDwj7l3x2hh46AlKxS5EftsQ4jTwTP+ojn44EBSM0p+OVSX12BKUvY9fU7+wf+0Kz1q
aw3Ae/DbnBc6Q5/ijqCXpVsxoADwTvbkULxexScCxPd2fk8bIomxQXumNG0ZzyOme4J/NYlkpgaI
qe9gaJslJIlhm0L+RrGPEMZ4agnqkhYLrS3H0T9yPjV2+I5xHVD0Wk3xHTLU6DKQa/OAAypoytmb
c9c3ouFRoOs0kIuLH1WxsyhNXObecNeOheWVFdpQooKxulyFvanFWDaierVNCPWCKxR21Kmvy1bP
6fMSE1yjkpzqv7c0oHinPZcQGjKGAX+SUIKi+sz2YCA7k4rqLmWrIQox6kRf2Lxl8BBeupjfHm/C
st0TbCiHt35JlLmlXrrWmAeo4f1hgabCwIgvAA+c2EZljw8JuPlCFDM04jRK4ksRJ+HrFxNitEfQ
44WjNSqR8Ti8MeLQ/Fgxiu6BviLB7Nzo/YaWEMcW5LGPo46c/TilQrtMjUpfv5/pdhDH6qHSK5RA
vY7fhf34CPI6mMiCufwC1XaJQHtSIImAwPAdbAAWyO7E4ivkOwBBddvyNVEAdlWu9foKWP6Xt5at
kaEKPGvZAhsK1J2wS4SLpMzAAfLlKWVIQiEhuy/Wtm9rnj1gpARHLVoCb6ER2y28csLD4RjHCjsf
80jVLOJFtxAKMdDeHpmzCctb0BDhLcpYlqjFDxkisKU9ABhT9j/yfA46FAdwccWX+3LfcE7LUqWI
GPnsglQppgoqtAjwyg4ewbUm6S5OwMtzAz4gYFITyF7HcnkT/7c2/E3oTLcds7qYXJgUy+X+Py0h
TB6uIeMWrE1dshriSqVNLy6rjY9cgAiffbwcggPShipRxjQS8054PL/eZdwFHoXtvdCd+33aQQ0w
zXGvkYT0xUqhRnel6CwBkoqN9mvrLLHkZpUDXyAVAcc1+JrkCpcoY3bxhJgMD6TBECcRq0UrmJOF
H+7eCNzx7q+r1xd1QGV9YlA+WTqqXW+ReMSq98CkJjWENmrb/856YLNw9vIOvOJkrXdLrIHV5bT7
c09jKhxuwyIHmu/9HtOLPe92G0jy6WV6GWdiYPmsqmn3b43voEkEMX9yD28OjA13bFe94XVbSHCi
K95/mq5zjjT2Vi3bsV95g3Zcuntea1c28bVa+ju5zso2poEIszicenkalyFOTpxFPSuA05ij3u8T
D0dRBhyxNcFmZIlbpT4OBhUIVQRhSjK6/FmCse4Fzh29h3AUqie4yKWq362wWusgnl7Gvtkx7MSN
l/E+yKrv2dRtcRRtuJ8qMvtSFCdDdtzeMPtcY6Ki1mg9nKTxhrdenpBIFwaHaYfNYGJs1JDQ+Z04
pH0730M/sUXcIsAQt1Al8Jxqa0BsOJw9jSfroGYRQuYliACeWmCjYWluRh+V6gxEe5+44DNOd0eD
XX60o+xipuDkhSsIv7Lz+GiHfPUcXQS8yiPz4wG6XlGdRbAcap8DvPTulFrt1kAiHrlnilGRSWd/
Ekn1gKs0qiI3z0uHlkLXXaPOCjSvw3Lu0dBIXQu2N+7Rv9aPb/S3JNUY384Mt5BT3mvkSsUY+8Is
dMI4QMCkkAA1MfMrOw8MJr4vlTdAL/4WFC2B7qft7wV4QVFD+f0DB9cb7fyAq366S20ovXywywHB
1K2iglApRiZFof0hPAyS+NgZVrVlQyJJ9jssiuGsb/pN+QH9/sVjqNabYNtGpqjmdJMh624cA7cr
PVdzr58feQt1JNp+zBYdc9zNHnLvxxFKD6e2A+d1w/008PgR2DcpKD/QUiU3vS8B6+ZcTs1zey+C
nkZrNCskxN6bN3GvBh/tzu4LckuF6uEm2vcr/ZPvg7Kj1Q/egPAdeLAinCZ+daxzS333X06I2fwy
W7YQTKRbSpj1w0ahK27jA/q285RQUzKJiR1AII/8wrHy6zfhmB/o2hnEKbt6Xu0UpjML8Q6b07TI
2CLGuZ4hSzYI+RtwmGIsNHZoTtZqm1pJ3WWa7b8mXaYjwLJTFdXD9cpgxsqQTOBs4Qt07r8liPmY
y/HfLZPSdTAO2P0Z/+xrD62n2eBoC1n42LurpFNFuGUg9elhnTUTIEl6wjKA0ym8xejBbSOsVn3v
AP3CuVZwlB816wIvUy2cq1rHvM3vQZm8WKoMRYbm992zCy0i6tnUPO67KVvDx9mjEUyru6WmPx9s
Ul4C57Z8i19CfEnlbQVMMhjcUujHvyo5F4Bi4IUvaB+jY5fTJlQ5Ez08GTOHVPmzxTnZUDlSbt8J
ADDvx3W+cGfWmaxleE1fGQ5CcBWaTpftOIAIsk75qWHbwJseMOeitMZRxFleyd6QYTpPmJS0KX/T
XgVXa/iyrr53qkS+gCIwLccP2Y2RZCH15lucvK8BB7iJCr684AOJjR4osHZtnbaNq6bdC86hjXOC
jicqSHcTZbeWRoyY3QOUGRkElMRt0VofyORmnZm4sXpsK3eQ1gBXOAD9JvKPcZhb1DLgRKTa8jOB
337UNzMXt9wEEUiC1m4AHkiLVzW3b3LdtWAvD38ETJmnOtwvrVz/BcwYBPTVEVzBnDF6QalcuiUu
0Xe6vgF1r6s8YzV0E81YhfyevzonxZgnw85fl5U8C15h0YpftWFLdttR2YnJIs7/CdeVwyB7dkKa
ShkUV3wpAxZTM+Ow0tMQOW+ovMa3RDOI7RCGMF6zuqxPLNfGkx5pyTXFxn2J4hPL/PKdUGv2q5fi
Thp/wpia5ueB90PygB0xpmCjoeHjnQb4sDIHwV8vtD1DRUsk/VerSYWy6nruPZoewLTX6PNyPmOZ
RwD+gY5gWIM1NZ39A57AJvCBNPyWw0MsZF7nkKEMZu2lRC6jB/kR/yCL/9FrhnI7j515dEmm2A6o
b5xKfiqYhLL1Td+tf0V78+x5LRmJImh7wpZDuJwjEL2cFucr/iBE04hy6Ha/dNOcsPS2ya41Mu0/
aY+VzB6qPDY9EhSvATS/nSoJ/9arAYomx9rTtie5SdUJAnHyFux84zIcy970JzeskDLUO6IGt0jX
ZNERvKZj99PdkyQGVjteNzAaPfTRIqOhcAn9/F5guzxKSW/i6N7p8ekfGv/6u0yxJIacdAEl3Okk
uM2eEFjkBr2BCJznfGF0+HyR5ypI2lHS8NetniI8SJuEK1EzCUl2MaIQwQXE3og5wyMakAoC7/Ex
ImUknJfe3RweLI2+829+bne6I75VLCwHcnInvm/BUGpVbPHEVJpgzXEVX8IhlUrv/hRqujsbFP5U
nj1e+JcamRnOqlHc7qcfJoFUMFfFKE0CUnTIoCICXkkrEYcpDbdcX4MNxGDFBFH8uc6qiQYPKQKF
tsGWvVgNqUecvWXvqpON5hypeLY3xrNVHXA/e0SODP9XT7zMCWPYQHX3KlEIp5B5aJ8xFUQzqpEB
OHtLPL3itlWQW57uMbb5y8gjQhwd7S/ovrT/p0frTs54laiMBUVtTQlz31Du9j905NPi7t4AOXIb
gwqpyFgtg35huixOFiNefVws6G75NmcwIKTuKMNVmVDebAzl75tCKICqtIb0hPNYkGDgJuec5sXD
jcqhvLXrTTgkpEuGwO+UKrN0AWu2QZo9f5DimdUQESj/sPv/jpCZzqsFTidYarsPte1oP0ekKweA
U7vs8slNahvICPyp80K7PaLsGYEsLxxMxdm9ld+6p8bzISGO8p0aTXyXzr3lBZ4ssH0f/xTfbAhv
9wuSMLDQwpo4hD1+Zo2+4Hb02ACWR8ambfr2wnOC0RFgGDGdm0PZjXbnVRnj2I0jlWqYXf+QQgjJ
I5Ifdy6MzXYJGtYbB+LR/byE8g92/d3ed9Xcd5LYVTh4cjc/Rw/dFwQ51KyACmKRlnttPt28wMoS
sn3DFVZk2pZ+mHoFj7DThVxNK49OCIkDp10Fm2LdxBCqVkwqnJvOQ1QhisSmv0yMGJ9Q329bCNzL
toVmxNsLBAK9uiSYa4WT6h0QnY4o3l0CTdIMXPcbnoOjewzhiYgvh2fv+p63x6Cg/TCvd+FfkGuR
+4OSdKkZTkOMfVrN417BPlBX/RITLMK3vmgnN5zeWoSgsne2UmyWkksuEygdPFCM0pNBkJ9aNrZO
btuBpq4tdUpVypH+gQD49AJVvrFrd+/N4XUvnFgvTSAhEJG3RGXnLuVab4GPmnwJ9lcAiN5Cdb3G
PKvgvRu41KAkeDQ4KQnNg8sCowVubjK7l8jkCLhwpbEfzL76sldlYmCjFtfB67YwrHt0K3I1ovHf
gWF4LlKzjSUsk55ZUtqwe6HOg/+9Xlw6iDrvrQMkRsP4mnts/iNtgjqHfNZ5uWHT1qoCk+bNvFAh
cfuxGrC1FtReWc8OhkNGJ8cUx9kpVFpD1PP1akvFFTMQmni4rBPoRCmXeuOaupydg2eJ35SBlh4i
wNwaeF7WKtZsA9T3rgzshXoPtO1Jv0ooVnlxL4nAgpAKeBR9Xi1igwDZnjy80EWPxnXrNoo5IR1e
5Mb48s4FkHa1sw5GP1Mjahj1fbimYnINw7ZCO/H2ZpGMiao1R51yRcpqu64PcD8ZbLaQMpowrWH9
0VgVeS6pSb3NRLat3lYDyHUrmS2qvEhlod0yZFnlJEgiZjr4w4GATy4x2ThJvxsCr3GT4XRkKMql
cvUyEXE8gz6Cc8KtaecPnd9kI2X1DmrQhepE/GJT4Sq+Rg3KwL116HuSJv7+IaAEaFa+IS9NCKwz
OfpFOPPFCy/gRSm/3MABVyFD7EjsteHEmXNuDQcFlnWRgIOWbjiuLluHIu9h+izlY7ovMaK3kGjD
2JC9Qx7WZzrlGk1zkd+kvmBoghilGhfa68jdHQpV0W2FXF0HrvcOVy8u+CNLDEnabJJQ+vGGtjsy
3FrIm1uSRLRN1y5uUlz/jlkfEuQiBjIbI9YGaCM2Y7iM3cDUi64vk5nKkiJ1iAdS0TxSbZYnJc9G
7QW5Z0QY8qtQLAqv3RCTSFmAWq0V3+0QegwRwio75IviDyfmitqRZTiWhib2aYqWRBP3jjG0gKZ5
/lzNEp77+eGcrKvNxP2odI/lIw8W4I00ZM2Xm4Xga3APOCRGRiH5MXHFe/HvIm2aiDVGv3W9B6zF
NfFYUOrDOjJaMCrENUAHl/9FK91u4iIsMpA2I39RYa/XuQV8z0Zy73XMkfZEoL2ReH+1uZUJdPQ3
VcTkE+QvpPFXakliq62u5wECSzXh0ioISZJTK/qIVZBGpKNskFq+qa35CNTWsDvjSDEnPSqh+ltO
tg8ukXircd9Aysp3go2W2ozPnTm6cCbWNJmf3eVEHVzVMKV6z81PvKcjZvVNpuoOuEDWFIpMEaX7
8x5CePTtFdZuJbJxQTzeuY0biQkHTBWqtC4Tkz873HLc7iMgTDcQ08u/Y243p4GOKAqDFBPyHhML
1zelrYuEy9evh2xv7nRQuMnLattPwAkqeS6dGu8urRnl6dUU3GLgY5dBOpVnhMW3zf1N518Arfa9
j0VxLxoOS+gKf/reU5O+ZXNRp47HLaoIrpSJ6wC4JRAff34GBrNLUe5acmcJq4dAe2bsPk3lPyg0
mqwEk5p+f6tzU9By9NKuwtc96qDMJAWnGtpMXVkrmDSzbDl1C2apt0gSTehWk2V0Tm3qe7wI8Kcn
i6lZ0/pzw+Usu0/nvotk88G1gpNaNXINOgmXPW6EGkoAt1S84MJCaxJS6ga8GSZmBn7/uiwYeKpW
ezbPG8Ln5guJfvPDV7MMhltYbTivb4JFyB3bgAIeeTMJUa9TlYJbskN6EKCP6bRUQMVT2CUah/rv
22cHgG+0DDBcup8dd3Vj3M9dL0P9IVHar1GlZKETv8wgoK84blwYf8Lc6HEiqqBSrTrFNrZC8YzR
uJKb+kzU2e9kpk6+6CKACVvqHf8VaWXzzsMrN8e4+m0oC8eHEzAnvgMzwAPEOW9VqgSrP9oFlGzV
LRK+TvMaWMV8i2vRSjXWDVMyEwdOMOGEtkzHaUK0TFLHgYBk3vJmQo8PgTmQpCEMhCfPsb/gWT9N
K+A0PE8k7vaR8p/ttCf1gGtkgEP79eP7HyjcgHflRVYM13EDLCvdiV8Sl/9CEayhw69/T7mlXkR+
A6tt1+ql2f6PAxcs+twt8JvvU/DVeLUJAVHc07IhWNjOlYZ4qumFEM0ssMXrUMSUxQ0Vc2Ft7ZmR
o6a59Cy3TGmo055NMu5NjjIkEsjk3UI+OU+atagBGc7sc+qGgGZg/ETRMZNytAf0AXszheH4lYxd
Q4SSrvVNesDDM6hWw3lT5YnybcYApGwYds7+V4V/kF26HT3xYtQEQqTa2glVoZ5PdwYyKIQFNNcO
m4Q/dxjPcvfOhbWp+YybwZSK+bDJKpFpiiYrgH4QLgMXZ49wir9DBzNgn5eBzHXhLu+pxnu9WF1O
HmyNVrB5gB9ko6ibWgpqkuSXdhVMINTWKFk3sTPaXBCAIf3owAciARh2kG8ww3KtMMoxQdjRTBdT
A3u/cM29cM6qWjH0eNfJjdN1flVuPnzpyYUC25Apx9z9ujihL3w29hOqT9wWOZNjo9c72iMQ+Epz
vTUd6rN3qxXl6jiIW+vG+kucZKLyQ9XNs4k1oFr1rkf2VjpZvLXhd5Lzsr4tna+vOOGMG0Q2pAqI
1EAWL9f6jH6l8Xb/nIyJzrBdLDn3O7eTXGYM9WDXI6oAaDpVVHdDzOLaDrufEk8uy42jnDNKg/h6
Cc53nCVVlCwTiH1nj+pwwPLgC1ZQkB8QjNQDe/kTWiuWsBqgz0I/F3vgIHLlKGpI3y3Kv1F/1Lpw
ImhcTcJ7azmsWm/C7+2NKhXQSsO78VHJXC+VtRX2hgnYejQB2QmrVZsSdNVmhAhzDFud4uFWDi+c
M444uxVe9t9FM/gW517n9ZbwoSe4vzQcqbYlsreyTXSVYOO8SrbmUCQQ7fP6s7D63FhLN1O1KkXc
vajEsybyZU+evrQPugBYCa4xQP4JuhuNjVHqr1OR66Q4eCR3c/JOtOqYw9PAVRMNcX7bL/mShQno
QRtDEh8vmX9KRGMe7DkTooFpXzLYviez2u0+kp8Sy+NDleDY1cibTDAP0YKJ8G6+vnjzjWOjNiRc
wayY895yHx9voYhkG+CCZObUOSRmDDzkwvB4nNN+Xg1TB6ImboFPLTpMxk2u1sMf/IojQU91SRen
pM8KxtZ1tvGRlMZjk6ftkiWEnXlzZRPQYQorBX1W3vMBGitt2n6UnZHBdZBU/7Ets/6oLOEKeL47
qSky/ca1TklSXEAFczVxLElQlB8gVI2SYFCoP++qxQA66CkNWam+L8aZm0km/o8NySk9rHbpK9w/
20Vr1uEFylgZvtqpdO3DDPVdSJqae03i8ihCxkl8MsTD8WP1UIZRGGiFVIHN5MgqE9TrWA6MlQNq
qfdm6ni8zJsVD7KIAKZZ5bjsYXONYCjypbpPRQfiTdkIvULPn1jhz/w3CMLcGBf7qauu4tnIvWBG
to9MDrgRosegzjJuGEZu/tqAEzAWE7mekF5KylflJ5iWMaI88Qn4/HAcK35ncdRLKr3rUTbvJGP9
qehXr15qIzmUJCzeqpEadSxa/judp8Vy9FVJL1r0pHX6aPEx4uxarMZ6A0yuAuLTwwrwxqDhwzl3
1DFP1EETAmvYLLBVONldij4WiddzJ7Lt8xeoFsp98Mthy2K3/xuiv2Aw83F/VdSp9xr4WsG2IL7E
JLNLEtFF+zAPBhKAKzVxSy0Z89xRPUkV3rMNQp0DFZmpy2N5D+A3SVqfz40nI0pwFYlVw7dzwQ/0
WTTmLETfX4UCZFg5usXruyJ835WB9a6Y9kzxqpan+c29fba4/UgvZImJ4R1CsqRUEqa0MhvDL8es
JQ4tyR/I1CpVUcWLzCGD95yZ7QMCmvl3hP5I5oKOX/oGiAKqawFShEn6lzOihO2wObJF6wJ+34Ed
mlQSLB20yZoK+qf3rPCft0NNYPbrf0XFMtNiuT0ax3q2XpGdZxKZrDjH6MeNDXzM/bw+LzJHzBwZ
ey7kmsfRsveXCMy0fiv7TZOND+Q5SLxBKPeuisdrsvYuMEshoYW85Dh5Meily6hFHQ9Bz3OocZUU
OqFYPwsAvcVOZMYJJIQXEehRj/ZgovluDTsIuGVUqvSxG5ifBUD37AdeoqYK7dufAzME/AeD+JNt
oqOVmbAFM2wYJClv1gL9kDCTM74F7Nz5OEiwoMGwwqiWO5SIGbnOgHV9ZfVrpaoUz905NHdptFSQ
MqgPnQcqxEpnv1xyQ5hw2YmMo7oJx8ri5hh3EuViVQeuHTtMGxrcIQmWierWs+BnGcWupyfVxfC+
dbrwFXrDi++EpZsE8JFSA+QEDJs3Oagm3yXzTuyTF6KON/l1aMN9X4XTPFdgf8qwN2DG+njT6cxi
2Q4mK24bifmpWqTtPe5zB1et7U9dAV7+44vR14Pif91ED7kDRNeJOXtd0G+ijdd9nP0XtgXPAHK9
NgEQOfXLbnoHYFiF8eE+W5G1cdHn29kXtpOBT6AWeA57/M4QRVsYktKnE30fZVuHHssHZKhETNdH
EMtEXkvP0NYMN8P0isXVenKCD9BtlyfgHWi+P8Kef9/Ks5clKxYKOhpLoLgRD1U983X49Ld/yCaO
M3XUmiZzWLBGuxbqHMoCUshWfQwlhoIHvoEd/LMeU166NxOzxzJ+qwC2lHA76jH2r8z6SpPcvCVj
eBISUzMSYwC09vFzmPKZCVtIkHYK4laSguR+5rHIeIV7/ivm7slSfQTq4w0jzcC81hB5u1R0UvRh
Iv9PbkLuRreruwtmKvB6yVdN6Ql40i+6hzpqbORdyS+7ki3LMBBltsKDrNGw9NxmToEdwLhO5zHP
ZSFmSDwZSu4lXUsiR987UOGI70nNSLTLbqsncd49ghadDy1BWqAphi0Iy5EBMQuqvrqEn3BoFuWa
CR+LdqNaLkw93Dpy6yCmxs319/PdYIIRwBkAmz4AG5fDAEI0uIOsWu4oHWGOccXjKDG/Fug0fLqv
qLIVjMe6XxrFeAvEaGNNDhVD2pNPRf1oAZRi9iwODyjdhjm6WOcuM/6semk8enW+nYkoLTVe3s2z
FMQcGjGIdchnn5TKKEavJkIAIKT9Z2N0NuSZiH0niSVnUGU/c+WnwDnhXzTUnhpR7254BI8LxgMY
cblRa2eBO0dhsfYIMUcJuCPrW99SEdE8Km536vfq1xInSCg4TQfnKPsvkYBA3fiz+WDlZUpQSgEi
EKCUP/iuDcCd4qwAjnmJqLDoV8MRkm9kRBikPcKfHxEOARJLxMPA+bIW9oOYHcpGGCIpTWpBqUdd
75/WOW3lFWWTXv5FA3QbV9nCQd9HmnfK83XvV/HFasGGg9h+N8+HgEg0mG+H850zb83N2yJS7AOz
RaOWYRnbvZ2x2BVpMNwNOMzMlMHfdg0zjMu1sp06PY3t4REx/c8jL5a59mdoBAGiB/rog/Me6Spj
IVHsW4+K8+CGFKfGb8UzecJ4MUY1GOOBEqFfniCktyleuCLRukCV/rrujxR05JaH2MDdUGWykvhz
j/5+NpLiLKxpYOuLY/K3PTJ/4ZF4DbcVHH0Zrg9Sjn9la0zGE7nC+rJ/C2aJs4dIUOdS3T5Br+Rn
2b7yzCMwpouA8dfFWRlppB13YHLfr3Z/VBVw93FTX7AhbN48V24gWrHLIcV+Qr4lPEF+eG+gzS3u
zX+LDmaiMupohtOCT2km6BS2ClvzuXKj2d8wXS2xBCmCLTe1/lLYMMJpTBj97me6dUd6l1LZESSm
OdmY96np09Xqx6Onn6CVNCxjGpo4kl9GPxxEBVdpuQDntsKaZ4BeTovhcM0rydXulbhDWpsqWdrb
MvyYYK4kmzi45g8j65OoOBEHsRFh6ym3ILr1F+g/l//7jUVthX4UIlVRuMBkAq9EyKYEu2c88UkG
aDUtF9koiH5nzHP7Xqo7Zz/zfMJLHsl72M7n8Ry15W2f5QxPEQzPdo1LRrs/yFLSPtx3YKR14r8X
QeGogLS27qVUM610sR9mHOYu32BenSUgxAtZ+Kd83pEmL8YudfTfYgcAVhtm9Br4KX9+TkkEy+Sy
hF4BO4vbyu9WLh21gEf7suFqebROEw8vqDAI3KBey1mejlQQvQG9YOXIQYVIbkGR12uA5MxYFLWg
6bnbqorseuNeFqZ/7NXFN+OEXgYvZ0mfRjHpUT8ZxYF/ACh3Bx8tqLTl44hgdAV7SrVz1hnS5cUz
KvKuC6pUWm/OhbFjDLCnEDFov+KT0In2HtTe3VNm3Ll0GgXjMctcxdWbNbst0xXstLd73wpHxBlG
3UIHpV+/gRIyBLc6wDUDrJ31rn4yQDQPsKWjPnTxfoprF9xyVWeuahUxzsJUcoFiMCM3cQvsDBfn
1vwo1ZpJlHbRQ42jg7bPvGnTZabNQdUMHL0SHvywFwHwh3vDQe9SgnTPnGSJjesnpcSbBWGtWy3M
7hKyxXPAOF1QKPKM1TxUxeiddMVMhT+LkE7InB55Pup2WstXpLblu3PyX3oZ5kuiND1YFY21ol+I
BtujgqEScghd98JKKIs02UhhGVSnALAJBVd9HWfk0ti+gBq81Ic42/K/LQKjlttDZ3/HZ9IwEdmA
RwcAdz6dTlTZiTX58MoSZNcZiCOVSKBTU2XmPToD1/uMZBJsvplxJo4j7rkjAF17+bwXVcJWvbu6
bBYdQ1vjEL0d2dzdN7vt6Mugs9kaDLjrmLDXYrjfZeWooU3iiC4nqJSU4NcAC5uTtGcBSPbQX/h8
SUjf/JapXnBSIh4sPnR6TpFR2cS4oAYeJbp9f5BgMoUymVtnvMC4ZjsuQ4mT1oXGaFh+dY+lwPY0
VwHoRnZFtJ2q2ZYSWOXUn46R5KA0azNy2EAij/RgLT8wKVvtjRbqqsCs2uFzOr0TAtyd4D9UVO/y
Am6+abFwA1vszH3wKbMd/XPW8daGGL6+UGyq4Y5tnsnSJOa5Z89eAMW6SnAp0/vOOGnn/fnXFHoa
BZ0dcw4RIbD+7mlRK/E86oByZAkYbRARhtTAprmwuSlhNPJaoZZmkxqCstC1gMOHN72sXZUkq784
WjgSveeIdAhATT0VUjaZi01hIZ+gDGg5Sm6D2wN/NHSOEY9ygp/CH4ybVD7LH+XfWJWLTxtmOXWC
HYuOvFmFJEEEuqS2mtC1xnp6UC3UCW4t+VndES502vk1cMFpv2GRute01cXweAcEZqVQdAIp5Riu
eaEIZzzej9FEtqoCO1th3ykblfA+GHDGD1RWVpEMOnS6E/jhwvwN4H8DlFL1l7tICVxGf+LhB1CZ
kPKi22G8NnjaJLRS0JtZ+qvnQM06q3fwWaUg7eQbK5PrsETZdLRxvvUmpE+BzUYbGUOWR2NtMdX6
7VuzDtStpi6b7pfT1wNxolFDn4OpdSZXJyavtYVIcBc9+RS2sDt2oWKf3rKMtxkghOwpkhnvtgUO
MrqrXifHS1ohacemMKAwKChgsJSrYk7ka/tbj/vP0Iil01sOV/gm61K11fX9p111idC6Xj+lJVIg
U+Vugp0ww/j5OynW05whtwHBRiZa7d4cHYvIJ7UcDtRgYWVAGzBL3p0M4/n4IAXVvcaQgSp8lFA0
DxbI8sDG1AaUI4H3qT30Lvg9vjYrZyA1EMBrEavORKfYQHKU/W+kOenEwC5gbwYRWqlySSRpNHi0
WuhyS59SgsnNzIZRaoTzbBao3z6+IUXn41YqPaKbJWQ97LXdOcwh9jU1IkPmejbrRlnPwZnRNs5X
x73Stnt+wtE8HcR7TKeH3lzhLgV3PLuPiELz+AsjCKhuI3ncYegdhWuosNH0okpWfayAQ9e2K341
oaKzMeKFTQ0bxB2Nw7UXlPImEHDBJXY+anqtRF2iMANnP2SHCIrjqEk6KJUReTcNAHqQ2VsKlTCr
N3DCqNfLpW5JG0uDug3YSDP3RBxLppvQNY3KWU+8AZ0kos1GVg7ppTKe4Tezqp5XfJWzZdB2An71
RvpnnVTGOrTqnjg/gkDcLX8dkREpPQqWYFnWdsRHIYQVGHO8oDYsiSdyUu7aUh135tVUK2xLAUNU
Jq2DKFeixFl0Uw8kVA3oHMTNjRgHt6/DMV+WKfJUudMLPGDi2p9kZbDtJvYLJmHn/jEGe4CPD1lE
m4dc4jkI/O37NLTmvnvf+slU7qI9Z3kxsXP9P7f/ofwH6eCKvP+dBWy34LmGonMfhceaYc5N4p1X
HmSsceHrsVwt0Pqh1MqQ2LBbHlezpc9lceDnDE8E9XsDEW/2raRWGXjIkCyCY7L9TiF6zG1j/iFq
XUMWT5KXznq5rITXyj+GnUDcLunSxO5v4CJxNakhvtCZtXsJUELsg9Sf/c+FdcUaadUwC47NlkSG
BBd54g5xEDJOF2OIDS5FQGnOfhHhOa1PI+HtcENWQVS03JTvjybhP5OaV7YwcovXFjWLhaNy6+LC
MzaJ0YN8V8SuWgzCLbdk9CwSZVKBgA4JqbyagbNNH0jlp8IdWhb57XrfEQxHs0eNsf89cToae9r+
+XWwn51PDKppHvFOuEX+esREmFwj/GGOD9Xx2T/h72AtBXjFc2MY53Gau1c3omB0whRjNzS+4gKi
avmtpOV+q3SUkkTGHf6JiRwExBFkYpWIGxnuD3bUmJ7XzAp8XS+bvDvVhphns6B0nYKcthFPZ11p
BrryN/DNsffV3rz5Iko6V4fR74voTqQS1GScYGwdlka0kSEAeV7BwIUAioFYV7Gu8bDcmWa+lKTz
/HxViDTnGVfNVi5mXlDsUTLAkEnDjDbhcAgMcSPlSiPuRgVdZWSuq2VIwVvsG90E+Y75keCKLMRa
ow0HBPdtR4sdmA/ua5keNK2gmgZvH+fruV/d/ziBbOJSM2EnTmYwE/x1VvbXQuQyCwNmct+hAfq4
8KxQO6taaHrqFS/WcmKEYPorCIWPPZWKafYC9onXKog3fU6ts95sSj2PJZ4USazXu8XDMwkQjnU0
ayMN/4MpfaTleaBVn90ik/hy6epwxv/27t91peDQpyvPW0JEMZVkVyEmL2Z9Iy8bkdhlx/aS92J3
5TzNsKgagfU86JMpmyiEPwXNQn/eRpNSEy9HoMaG1+YoAlbCZac13KQE/xevTw/SU4lbJ/baCds8
cD5viJSVkg7EREvyEaGXBtcNGb9oVvqTzKl6I+JLkTF8FVfSvXaP7nAAbUek0tUob+jrbWSr1KOj
7v4ZBKENcN7VYeGZXcbDGoaSc0rBDME9XBSDekTN2QviGX3JxaUZUsSsWyqWEtG/F3JJ/QFMoXkp
SoUSa4FXHZblxwapS9BFboNrJj8PPlUkvHevU6wklPPdpMPKE9ZChfK1F+kl1E6q8UIFUvhrs+O+
8ojude6BUaMXCHELpW0jWloG+uFbN2ZuDcE35vBpF6ZjgR3uepl5EcIQP06/Js4ca9M9ixzuV8I+
OCGsyxE+mBoFdi8svVtmBqpHOGw77JH2h6IBjDXnLjFiYtNBem7Geh+vufdjgWRXURMAlP2k6txd
x2USq9vhQBNLWGtQVoKQG1uHh36Jp+Smke4csZgduUSDfJGf/I2aTZAN+UNPiZkNKVPU4XEhWDDK
xEXWYvfvKnG5oAnx0oQVgx+ykfPgzV0XT0Go6JsinJ+Ew9RLa/o8oQBAtoMlIhHdX+sco6nFU5BW
l6h5cLJnYCx8Wpj0dMUxx0/JU378ttFdSohYYdXHw8Q2H9XwobH+C4vSsPTQZmsq9FK+xSFicMVS
9BWj5hdMPnRJMC3WT2mxNBim8d3ufScgXj3ElBT2nUV6VeIHpi3SAG+kjxouVbUyhadDlyTgO/4w
Almm9hf4guxf8pORWDAwYEQy+K9VqNyUZS9I20Gt5Bk3v5rzDTV08izbL6otSWmzowsg+ulY+FfF
JmPALxOSMc2bN7j5WHpK0eFBlIKnRAxFTsFgbfBtEwErw2r+3Cufpx8I3FKfvF6i2W7CNYIZ0muH
qDi+DWCkpULDjxbwa7aTjAii819qWNbooLTSecqw6ruMaVCatdrBChCM2JTgj3wQgumJg5mlNt8s
DD9euTIbHDBPQidN1WFR/gS/AwvSfIBHawNM7PJxQx1JseVn0VAOkJYd5Sd/dTyqT9wStHzMTBHJ
G/3A/Ge48nwW/7gWGl9+pfQHPN8Mc/D08r/6aXhXHb7KbPqxy7Iw3b4QUBbm49zVk1+QLd7/1TTs
EjKk3jGVKZ7+bPHd4UBAs2ys19pZ2AQXphmPNV1YqviVfxIYuGkKG8Mq32c7SM+kI8qu9aj47669
VmQCcR1oNyDgaU3wRU0sd2YGegRBmM9PSAvt5C+mgFqhKdRaGUdm161gFkAkpqZjMnn7Ys1ha4M5
miwbLUR3swW68caGX2274V8cLIjsUsbDhEMMxJF7aInZkfvioHYmEa+LrYxDhDe+8f7OPQMSjc1v
a5gZPuYm8FXwtimsm798ZnNFpi6ovglrkv8dU8ZUqZ2d77Xdru90uU4Vy35jitN2AD1mZxf/MRcI
bJjXqL7MK7LzS+ElQ/nC8bX8xJ/wtHcPVOrfkhzD5krHj8M6s2tZd3HSTq4HYRoh702CJcFYRxCy
uykc+S3jg0SwnTB7TtNSS3I7UIkRixiTCQTvdFl9hGGqaRq6meg6eN/jHrq6f46AojPysvMMJlBG
XtAn55rd4pmCmiMMnVHyakIhrcLegK71IJ1y90mqnYAL5m5oFlF6FJRlfSgFDFq0oTMqULC5nFjW
IrCiR/I15b70XaxwADyX6MHsxOa3s/zTpAkduW4Fv2I5jFseCpwK9bgW7sV6LnseHpSuaEjLxblj
125fDXjUqskfAlDXS6oh3ar+Pg6FbTd/soeGxF6XYCSfEY0aq6cngql7kfJSrgdYzf1xl9O19NTc
OxkSksq/RcG4BbR2pRfCiZzqT6p7EJe581aQLiHqndMdOWdh2StwQDILIf3g+OwBuvzxn4ubZLFa
L5BYP4ee3kIjYRN3sn/p87e124KArU6uAD7NV2fO81rR6O1cc7io7rMOncM6osdlz/Ihw+KkeVdk
8mpBUpvsvvRGeLUw99M64EWY+j1hFkaVChD0LXYvRHKEwM7hM32rr8gJQ7ABVWv3ChPn/F+w5Eft
L2OV5R4pdIuU+TDVpnIswcqTBAMCeuK1wlGcPcL5gLQRMskxaSF+3DaR59mE94cl+RpoTekU55ke
iG+FRResuYjsAOtuJL9AEdwUgGW/EMobY82pBo8m3dDOLpoZ5tF5MyANlzHODQ/E5sE8W50e/0/G
2bPSG86tqF6ebgdBmkpTb+smQ9rWbu1t2Pvmf133SF84Szg5VUsAAbujKK/yDWvRebnbWAiVkBCO
ouhHX34XIE8fg++MP3RudBb7LGNlKWvwvQqD3Kw9cQeMUF0nD03SDYpdXGpPXHorEkYmLYEu/C9q
XHxSPGIkz3HmjL9q7581UdGqAUCSry7k/4WLepL1oKGWXNPs2grsiAaB4WSOua6JK+Saln5ZIUdH
T39jw22hQg912+raoxwrqmSGtOS2BPwbvBbrk9HXipizHLka0uFnxEkSEo25Q3m4FuluwEPQGhqr
zP3mIUFWmlKec5y6cmSuLFB9yYkqb7Qq33q1Ip81WYc0Uggpz5UWBl4a6W8NwmEjskTTGIs4sKJJ
c4YZDAvG5MlTmWE1J8fNgPsp4QgnnFQlcRUEy8XURaRH/Ysnz+EYDj5Vlse5c2jyARXpUlAizluN
4PZa3F9j2J7xEfqQOnkulEt1ZDubFX5qh9TgMmPGuY51dYpr1kStNibacRBCwpyD1ezX0sUqZWXG
7LGK3Ku4Thq4veftD03kQNoVPhB7YYnPA3AjnWi9DpXWSalBKRBlR0W7IQzS5izjxO/Hv2ENP/Rw
Ma2Ei90Y0ZMk6FknrBjL4KfYOgka3sQm6vawJwp2uDv07uBGhbXDc7yO2QJk5ybLAfB9/8Snfsmz
wZzZKmjghFQYVOTNgqqLTkmHT2MjmAqqW+ck0dzhxTL8B1aXZX2q1pKDc0fw1dXw7xTVWsHDjlLg
kYRdk5Hj67VwQY5mYaAOwRkFOJmhG6Cb+umH1JCFaIgboRaDlfE0gyaKAgUrMiVJ589G9b40TFdy
kHTk9z0VcX6kJYvCndfETXt+soBnKTbpQysHAA8/Ffjqpd0u8Cv6GagEXYocL2k8+rIZNnGx1fTy
+HWyxHPB+S3weJnrIR2cCe4zfjiRLaFR2PfKdW0exCTbfhKOdhndyKNlHSxXtZd356y5bY5eGOoG
oo70RPlPoE/FturljK/TD10Jj38mNZFkayH75iF7b4AHVxsBlNUk0JYfGsBtZyMJYPYnSb4T7r6W
MtOTHZnsOxXN8+omz9rOamiU/SYGT8pX07i2YLtBXLKdhjIuXog/ZLpYmiFrC3LdAwrnDmc/m9+U
EmHGGmd91AP/ZPom1r6YevcoEAb6z6YDhHKDKrqDRzzepTmsLCcccE1J4W8MuPix6i5TNzqXPk/h
2vsloP4LEjkaQPCY3NhHfn1zikGMBl2rRL66iMbt6y4g5YGt4tTCOVswmgIbCypkZ7YezbEDOMCj
+KzYf5sc7Wb5cenaS0FbxZ9R76UJzROi4El8e83J1yNUhKiY/5mv3bhixzefQ1XIn3m/jyG0unLV
fFvADf6kJVkUMTAOjyFhgpI/GLpmXBh6lefHLS1whI3CAn/x1x1okkvSkNTMGxMOrO6kkP2tWw73
XsUQjBdJCh9I4BioXxJJmocPa7Jgk05Vd/d/FGF1hongJNVhGJAo4p6VXldAMpap/JlL+Jd0EuBZ
3MqHJXwd6azfNSGB1TCgdNiJBsO16Unc87EmXJqyr+yf1Hps0DkrAT4AskjQ1yxxj2FeUQ66P5Xk
3/fq1uyuC8UgX3xq6KVSXYGbjuv42rcOw9nut5NemxFyYQhmYdoRYhS38t09ovKpDiSqrkF7AZLU
CuJT4s3UmkOxpCYv+RNrr1rD2GHO/wN+GDDQ/WiGucXHRx6gzXgar8iyJOlyBo4xaX61SubmJyTR
Y4CS5PvVDCQTkQNVw99pae51gVuawkcVykhJ4GBdd4qywD5TRZguibuwRoVRqLgyI7ysuOY3TZpl
fNe4TUna3gPsmG17Lg/gl4M1+65yv86qInEZarqB9zgqVJtpeLoVFuDWyb5lgRHuXb5UOOutQWvr
jCanG0P0zRqsEBvR9jNhZQcfWfX/CGSxkqc+dqNQgSt16GDwzck76zzMR7nXyLHJw3rbX7C9putc
BEHb/q+fwn2Kx1FHAY2/D2lITtkskGk+jFH/vVSIPLwk4L6buddypjVnusnYoZTFZc0uKNdxNafB
cq1J8nA+QdTjzVh90sRhKK4LiHs7E3XCKsZT3ux6y1eR4w0hAQPuWH0DG4mCpkcT8bcFHuwRUKQ2
hW2jtGmaXjr1XqDzuWxKSRX3PFw/n6Z4P44GpvsdoVKIAzv/Om0EUW67m6EakZwcUTwpVry9LLma
sJ+LVPCZ3TYJCwg/Yxqh+kzXJAP6KK6+AZ9lpykdqZIpBKnP5/5w8SJSChIYvID8cegvckQECGBz
u+nCy861XtaXiCiWgA974kCeRhjnTNyg37QGJb22yBajIvt6Vjklvmvm6Jn+qY/v+iZI6xyvoH1M
Pqe/dAFk0byR52LD852Avbs5axSK0gBQMeGb3P1/ArO7BP969tHfLS81T/i7gdjThatveRRYmJKQ
Idlpmr9f7sv2Zc7qYhcqXaQWb3uLuSRsDQ3+buauRKt8FlPZgLQ7pCI8LCf4gMZwt46ayXDoStw+
rd6l9pCBPzsStZGFZklyTxepAcigG/qudy9jiAX8ub0VXMiHGWBtVFIxILzBpkGC28dKLXvUzLlW
t2gKPEZMAW8Gbod0MzYlU7QkE11lZRgXn71prs9QmuPZ3Zo43Kysue5c6lVItELlp8yUmwJP4F6C
ACyZl4FY8txWMoS7rC6Y1I4x6YHZzpwAK8Coh04wT7kBMMBVB6l7hANUGjqJEeW2qVpUuN0YRBhx
5Zd+wU/0jxQ9aMguM7PRDK7l3n7373JQNnsMNWGCkCeq3lCv4e6dP+PgeKhJoCfdwSDYPf1Ay21V
1lrJWRiBjuqnDE+angDRCfm29tjS37VTweB/Wd4Q+ivYckAtjpYeNRUKVM75LymzuVf01W4JRzlZ
KjHiF/uoCJIWkTXOvXgFVh75uv8EP/IS8GpvZjrknaBlMikgBKy1ZldAM4P7IAVWtTlQI5CW4dlp
Z7zCGdeAyzjTCY6sqPTY6uwJUsWeWcfukf1UZ3du4t1mYq3J9xFEWkkGRLGquqiuy6jKbKSRwRZA
kaoG43b/LXR93EEpPGEQu0KEUIygPZqHj6f0AuFXnxgMAqTYAhuU4wKLwx+WWc8zycR9H8C48aMs
T/4DqYF00by/XNnkEYe65fPhLAp2WzGwnECFTxBix5m7VzhQcQDdio97I00vg6CdnprsBLrIJTF4
PA2ZQ3rTUyk7djMYFEekNhSEX9ojPFoaYLpP/cCZ0jttLlgprHcDNK896+vZGHNrDyTp42G71V34
PU5LhfHnuUZFK1rZqrCaHDJqOX3dyJ8dsVUMelL8onZ17pVnZwy1Ngvj7QD5nJEZVGlGXptL8rDh
K5fLO8CoZQ/Z0U3rRrIcCD//09Ts4A/iRsZm4VtXFf9c4HrtUygwSy+zc5wzZCga/U2urFkT5WL8
ntky3rQc7M8m+uCuCBcNM9mteD77b2Is+wJnsePA98yKOzK/gUnsjtdAj0usYlR3s0myWbdVIvO4
TAa+t8ycDS3KTgXpjYf6v/EvI3L9koemJPGdZf0Qtt0kwJsr0ayNAyFwQxzr//lPbq2Ttt/nkXww
ZiBXqaTunQ1pG7hUMCC3NqN+P4x6rbe4u7gYgA5OjWA2iMpTVGmOcLFKQrfnAnZKKBaYxZ4ukkAP
5kQBZ2TxwTmqOKrc0f4bRoi4hKhrHqklVweO7wyTwdspyqZJEgTF4u0p0lxrorVxvcK33YQWDBr3
98eU5+8eCwHvsV4YNHD1RH6mpTg1rO/P2y99SjjI8jVs6r3VRMEYWwbjOg5TybujJ2Q9CGDKfWbn
IqzlMjqhxXpV6Px+RfMICAHi6eURoR1FFM+iHgDSZ91M88xWYFHko2bMcRgzATh0kM/oX1x4mLey
gVeC4cvoKRHxPwLoHgXiE7UZTm50gk477EPb0oBax83JDYJZNzyEDPUAyxVF7X7ZRQvuLvv6AE3t
gkoEWyCTmgf0tILgqkK88ISprYw0lp9VbbVKQTdPciHrhZjEc7K8oTDqUBXT+FpfAa2+yuGbkC+r
+hATHplZ7unFDQ1Usjq399nbuVNGsK0+nPM8FEH8vtFMGwEvHO9yQAct5obUER9lpE0S6yUmkiOi
HTsXbicbDuMtum6gP5MTfwUTSzuO0GIxUfrsU98dIri5C3B9n2l7azpBmOtib9AM7BeBYe9oLGn8
jbRmh1mG6mkc6TQC6z9yfdNfIRISDKZkDwsHm/difZI3BpcsvIi4gZgqD6bGUlbfm4W9Igf+Eca/
j8f3PBg10FrgqRhCm3/T6T/MZjuWLuQGhusssDiEX0UJnoh1KYRwnMgLC8ytReaeiXix2Sq6WA0/
3AyeOVkVAAC9GFO5F5BEsFeW66oZKY+xWmrr6ecq5NwzkU0/u/SaXbrXGerhCiZK1idgZXDlEc7r
uZQnVbLKLtCCZRZJ1YWDWAcOthx0PB8Vh6FieHYAZHL3TgY8WWO2l6d0+IztlS7xAdm+yUtE+JYF
pQTQgxpvkW9tU6E5WQcaLv8GDH40Vn+dF3+Eq4u5bc7CDBPKj6H3nMaI3py0+/AYsTq43afJ53Vu
AwLmeAWzgW3s1T/quaN26hDke/8/mwEvPFar9EMNSPGzgiH8Eno5Hs8BT27OWEQfUETCFMuHbGec
TM8qIph9cb1z0zonHMr0dCZOHwHX5R0Z7mS2NHYFM3XghgOfQ9VSL1TXVFEUFJFwwAHsPDR5+Kn0
KS1Ldrlsi+wD9zcuXZOK1PrOf/PipLUbcNkoULtm09+3f7ma/CwhWeYuG7B1eHXfpFfyMZJXoF4e
bHWbElGhfxzuL0PeymyrW2+kDevt9LrLlPq9GQaeefAQ8PVsauv7xwlYfMkOHcHvVcJnnoWYKI1K
AD9zlXLq1s853OLbO7cXuG+LeFBsP2U5Ry+Pmup5FuQEc4RtacpGxlZhvnyja/1GtHoNavaBi5TG
Rkq8AacWjS6haHWwPl0V3k9dYieP4nhj8D+esuq1NlOF6Gt+Y7eVXhG2YF29x0Jb5XNnBCyJGxAi
sv8cR+9TQfX9MGVPXl9ze7Fn9OC+PyI9o7d8XqBISoWr2EIvrOtA9fBWOS9fG8c7+WDzmUBsNdyz
cTuZltKG1tE4rzz7vDLHNvEwx1UzAN9VC+WHK3a7HA5Km2j8wkyPB5SRsVIs9UH/vR47e+1MWYdJ
szUJqluWUtmn9eRsak7n07RKCLf3gyCprVmorRuE5X+CCbRVrGjyYeIp9JV9OPL/RLcE6OUDgKeP
LLjWPK7JzmOnrurpU0+CfR6XW+aoFWzwcBVhB2xZ/7kRcbmvM6FCXfyBTFsNASoNdekEUj5yTZQ5
59X6ReuOMJBwwcCmJQPMJqeQNU3S0dyTlQYXacmhb9ayWvP5YIWEkBykSJeMiWuWR30RfgNf9r6W
c64eCiVqeYlLgD/SRK/xDtvltvF2NKG1XM4zZqkbqBbDAlk9UGsmL6r+/DZodTPkhDr5jWPxkwUN
b3uvRLummjGk+C7CVl6V04fGMaR6pKh13G3SoC8kmFSiZOwFnJ3BJRO2NNixKrqLGjG+01arjkzy
+JV9kqI8R8T8JDoU0+FUsZE/dIh+uuMOY9MyEgpOgp8XMGotr+hCgMFi07mqWmv/scwi77/PrmBu
HNrvEhd89qpJCpRi0k7h55LXHe29fv5GS04/UrUkUMv+kfyqHZqpgJoaE+TdLwFXXOZlq35x4RTR
Yazq4VIu32/tcdLCV+yEbHWZQmjvQ6QYeB7VSlxAlLhjhN1ghi0rCIESXufZ03gVL2vUfMB+ZVdS
KqsmU+ritmtTSa1shgzEGGiOVNzvf8r+h1nzVlQsZ/9LWv8bL0ORRNnOpAouh6chZcFe9Z0XPpGF
SBhTt9b8SkRja7WRdGIMcyCfwrLC65/BBLZxahFUkBbKOlTTf7Qv5JYwLRobScY0Tv6tG8mfspJZ
IOc1KkVXMJUpdPreEKz1xhrFiHKiVRb7KZoRS8C/kUPTCuBW2Yr7B7bF8pwdvZFLfFRFvSwedoY1
sCHDr11FBCjiQqFIzuPIYF13EJgIwATnLLzz8vUXoOR0QmLCD+wiwsP/E/q8J5XWaJ2O1vkI8qmJ
DiLGsRcZIkxLYrpc9j9nqQpCuEnuIuhBGbYgQC12oUkznCWmvhvtgrGAwmP1TUt22+pHt1qQH0lO
uUX6vslavdcVHDscYPwDxVfqcFIqqkz5ev+bXnOTcgTsLvvebDRlyo36sQTbqLpF72J/7Dkn4ydV
KjoGAflG5QjBM8Ohqz90XnFUteiIVy61QRwfUSBP5a7G2houKR1uvn73MKQu7j2zUG38fdu3551s
mK2wPBz7ruQhNdy3bcWlOXVjj8DL/R4+R8qbl+/t5+OzClBhALjsPIJKypB9yGufegg5f4U7IlIa
ybWnXveHf33kVQbaZCzir4scO8gIryyKQEgLPLbwxqgoRR6zn6uDvxhsHdHwe2hswT7ahtAzdmgC
cQPyraWr8UMy/e2UaPylKJbFmqdewa5bikxGQa2lhaOL+UY3sMxwbjraBdxns7vOFGntmjR0gq5F
N9S1gx+ZtISnmOrSZM+wSrJ2FaykNDI8hAvcolN4kGPocYBaWpZt1otopmJd4DJq+g1VUXVol6aj
c+Dwk37XvTYANEUWn0zq6OPl2XOnalf8gk6Xzmt//XckA5KidsbhgbTa5iZDd5o1ai8wSqZPnVln
DKbrY5DXR47opw1CH8AWNf+ORu7EAxWXm7QN0NXe+cbJ13Co5i1ygpPU9+oOn0WEupG7kjsdH//B
WMGJ5hJ3Pq72mz/DpEkF89OKS8HKno9c8fomkLQ8Thq69Lsf7dOLOevBPpo5wVp2uftkjVH4ZSHO
YFHhoN6hvxk2+yBBhut1KTa+6InA204nggmT//5yK4LCOTJNo/AfiGjE50XLYNB+4I4+ZPbUFdjo
LZ6Zh7xkvL29RaAwcgVC3gu5MV3A4SGPkk0pjN4sh1sPrLywuhmYle3Chj1A6j6lB+kgRGHU6cWq
bRGAkqRta6WNOXlOH73Jf2VsTN/RuvM5cwJ54nCmEkxA2uShqd31NkwzSw8evFfukfXMdFQEkMkw
RYDjqM89nogLJBZ5yhtZuG+rSNh4P/NUXspGnNg8sthrT1CTnEGGm4eZzMImCONr0eJyxYxnhuZE
W8jbZN1k5YTG3A8wmM0ZLCEK6HDHCrNrsB/+v6q4e0KING/24fl9yjNBu/cItIzi4FJZWhuSp4t4
ti6nPfISMK62+XJ7F1xsNE9eqijgWXSIZBZnGp9L7ve3v6p0LMmAtNMtvZuQYC7s1s1PNh4+T1ko
q+lqrAL/nc5BoBSIxEX314BhLsrPIk0GfDZZP2XTUOFA21v4+EI8WXx4o9LA45D0BnFjNCSOWxMx
ypZoyTCof5eonbNF9IoZianz/o0y2GDVN5RgXm2Gp0MRf6FfcDaQ+I/NmR0oJfc3Rtghb2hUcTKa
yO1EIM7EEJPus9ix0akf4qhP7XzjGZUxLyLCMEBLjyn3HsGQSy7zq2keYQoepAeEYQRBbUaABJM5
CVRzpd3E++YZup38snJ2EomPNHB9kT5A8LbOYntCDj1jPuxWIg5/ePm4VdflAufh6RKpbTgqSX8V
UoLcmveb2dOZeeY/B/guocmgt0EMibQwp5ep5moWHxIzUMCPNBT+rGaIPUfJpV+IxcOJ4ek0c5wL
v0fM62YrNBQjIz8VbQnIPrbtuVPYMpwgn2xf+83eJGHGdmy/O9r/QyhPVmfavGDjUgAgAq7OYSOa
Xfgmkn0SIGyK4rOeKVusVn5UphJ7o7TIDot/MGDlQ4smMaaizBQm2gT2kKWJBSS/nUpsZqsYYW3H
+CEsccmVOTxWHCzPB0gF3BQtPmtK65nIWUE3pOGEdzQFzNKyqSrzya2+fPaIvVIFHWMUurhuPUT9
MPrPsnkr1/+Stexd3oJS8VHWQMXVtKnsIKXahQTXY5wgn/rx2qwuDD/o446LKEDD8YuNQAnOXT5E
sXze0UDUw6VN6XRr1Ln0bCih0I1ApIopsqevUS9UFDbAzobLEd3lCExKKZLFg6xKvAsMc9fTQyaI
zxNbT7wOVvXjmZOAeHDuC8JZPqQJhD5GfVeXDsfnLFIbtLikDOQ5TQ6bD2QbeMsc0adQU8e0XWke
fOi0HJ4l49MVruQnxnTsq5my1dF3cJt9D+QZfP11Dny5lT8oOfXLqz22+qCgLNT98yKI7Loxu47o
4DjZ1qsojPXc/vrQ0ksotDzcAH2VOimBut5yVC2Gb/EVAnOcqdposyVj2BvVKKuFAYfkOAmpu8WZ
vtcmNhlIgVMIsH95vImdUzr0yuvcMOnPyEZYjNBevsD+I3MWs4BXpfEcZ+tzDhurfBSFJGkc4ZBy
gdbYj8aIS8CN2QSuuBEhpW+DdnA794xg97ia92S5mlBMqUiYrQ0+dSm25irznY7K4K9e/shCFpmP
KSjUMCQoiXOIX1szmwnMuvm4aJXpb5pxCzMU2t89Z2P3NdagRt97j+uQfnrnkBKUZvkrwPlP3H40
mHhusNl9pR4APIKDx669znWPYaoS6Gb66w9Bv7zvZrEnaUZtW9ZF6JsxzJE0WKYUyKOIQDnsfy/3
lvJRGlLNF00I2S6y/kdFM3ZuPLPakxZTHgtUixYXwNxGhZZpQA4DdaGnlwZqlbCFS9ui1jcTBJAo
gXINfihrqI+uiZUxGCzNQw8CY7IVpMGGfEjavWG5/0STN1cbg5iVVyS9RKjvO2hiIdkb6vyY2EzL
Btwz6IPOY/mwNKDXAy9HcutReChqIcreM+q9ALZZD8HiqzFYdcxgydCCREZv6Bj2mNoGV1jJ4eYx
mBGbgX8F2Ib4AgW4+GTrniycxRDpWqSvWl/W9F87tFaC1ersR02UVJmjDDwFQo47wCX5+UtMYSfJ
EsOSr7ksXpYGbjjrT4Lp6zwxFfnPmKYxr6h4elJm27l3OXRSqZu4j6/cNfU9ZDFpW0UWHwtjR1Ev
3tBRiovN9gmMZvuWAMkM15R3e4G+n/pUxtgOWipW+J15Vo7iQT308dEI/YAPnPXIEipFjXX3uBU/
7HgRPuP5IcQUT322ia5IOPs/guO38kOfaIiGuV4mEaYfWeKyMeLX1cYdtyAsaXgexwWPQjGqTer5
siRIDEXrhUglctDuZieYqxUAYFyPwrZbYyTpiTiNQH4+iFcKDvLXGuz2GT5z2L6wrOoFbE+ImkGq
hi2C1gRgp9uFWNMhedrWZWuyVzIqxuCsDidYAMuX/GVBdVhOS5T8Fd7sgtAZEGkT3YHECaMtGiw1
0X3qCYsmnE8N8ZezH59IZxihcN6kCIHuXvKvMxdMv5HfYYTaS/SemxW4fJLMJictVNGVGSp8EHOC
nyvsxgRjky1EH4KfWi0gkqF8/wg5wZ8dipVMc79woUd+VkOrVTen90GTl0meNE+NW5vSVbPL1Jja
KaiSDGgl1K2HsmbNwsve5VvgS9zuPlBaobX7iuYzIalnHXXESK6bbOxzR7t6+da7xI+YWdxU4a26
eMkA+wwlpBBZ8rjPcVwNebLVZ8tg3+HwMsA9BRZnz7Ntl3HQYFZ67qNlf0DB75P6fWoAb69WzUBA
K+on8WjweIx1tXsfM+Q8J5yv1bxBwsqr0MeMvfOr03HU2oRg/7bVt1ituHKkE7W3Y8hSlupIOjPE
arUi178i0ifJgG3nIQGc5TgMK+DzTNBWI+lQSTT9Hwp0sk7B9RDWIiPjUZeR4Vv6oN1+Q2M08ZWD
j+Oj0M72Gjx/JrqfueThrjspGF489b7eGdrdSsgo7H/deii6XsZAq+Adl4mOf1ZZoq9zg4f10c1L
r+bw5HsuoVYj2LD24VsBITCJ6fq4e4Tdkb5o2+xWnC7R8PfbK5wDMH6ZyQ9sFHP1dMzZVZiMLOYO
86I63Ce9IQsx/R+jRhm5qCYXTTddp+xThLkyTMRcdYnqoq9q6YUmQtbPPzVLQmbEx2TFpAYjQjZo
uSx6FBm0k3JjhhHSCrjPoU8qFfGXC3T9zHuJRFdD9x6VYlppbPoAu3lznwZqb38q2AxSa7rA2dGz
EedJwOOHqBnqbUdcfmJGjrO+6J66c04j2u8JvAvQNIHghi5ixY5C7a+5u23cRmZdGuhPaborF3Sb
TQoO/Obbw0CQxaLwH8rJYOMoG+DI9b8JrG/CGLFxF6oMLNhb/bKCrPxTaNpZmsGD/Z1YPHEj2fUu
NjouXWLnQxPm6EJdwS2IC1z53kz3XKb+DmU/nzUGSN/xNkmggPt2z+tVEFgJkZA9zdl11myVdH+i
CloCMZzEoqRm37sSJD/5/5EVfG5HRUEW0xM6N+Xd4kFMPQMgK4+ArG31CKOEp6hEVm68uwNK/kEZ
MkTaRtJg6spmA6rXAXhat8S80h6++fthEaqcrVEF9usJT4KhL/KiSsX0geZt9bz/8CBe1pzXah6K
QCVMt0DB0+zB8n54zyQEIvMa6L0d5VTrnOzAVLWuEIkJlvdZDwsgTZivUOqcFlR2mX5il3s6wCRv
nGcg+XI3RQm9+dge1BTC9mt//JROq+/6siSGtJVFKvCzCCujT7j5BbECdZnAadZy+8cUbD/oQ8aB
AUoDHYlaBRug15om4xhOKHsACr0+El+bomJ4z0QgVTklU1kHTSY1EeNKlHSN/PNKoiOsdRLu+Bux
tTlv/6lar8DQjnuQL0d/7F8NffxukIIQQNmvcvEyU4xsmV2MSP1WZMCKIp2EVYNBc5tfUz3Dtdcm
XGsS3YOT1KbFU9yKCZcCHkMfxkDwgjjBqmES5YaIi2mpJL5A2xmjp/VxyV9ZFRwOFgN0EYQDzmRa
FYnsNTCauCa3i4sBbLxj45gzdDjwo2HoxfLhWbIRfsGzljEBMKwGtx9nLEj9zpPt5dNMtbYPnLuD
8/TIMr4ZtjUEA9Br4fvuEbiPmVOu5EAf/BvkM7HDmv3Pulhmm1jUz/QYXxpTmG5Xloq6ZDXcXFpU
B0vcuD0YgjgNrp3tn1/Y347lilBn74iGNflwk5E2ASkz1WbpdsPGtRt53JU7Wy3jY3tcFBmTH7pC
qr7YpNTdUnwJE18AB8KmToGCfeC/ferMh0E+/bPfdnbFR54qmbpzrErt30CV98KoxZ7SNf/uRt6G
c4sEQv1EPzT349+FoQc7pLisShCrIU0SYeIc6EtBlmttevDIGXGdRNFVPlRAF06YqH5TdqQdWd04
9bH8Qqsz6Z1RHSSZ1uZy3ep3ESgnVBqWV93hG1w3yeb21eXsPl+RdciaKcWFpO0UuhInYNAb4wuV
7QqiGFPQG2SstSwuAtt9ZQFIwJPuCzjBgbxK3sbsSI+L7uZTKgJHSe5JpxnmCsU/23AWyAfVvvLd
0UYnvUtgqKyzPkYZT2tqo4AHngnvPx19hLhVj6VkTXp/gXYhoUh9QG/dOwXuabKllEiZpFtvATG8
4W2qQjNHAgM5UEyhCD/PEAwQjnTZU/BMyDJ5p6CVsjq1QXVJTTXtM5py3fsZRvD6806Av+Gc/aIe
Pwe/kaWiZqCniZiW+nzbti9XzI1dzXIwdwp+Qy0r11u3Y770gHbWYjTVv2w4nxoPSwEjevzryDl6
dDT26ZjcAmFU0NrZUHGWX57/Irv7Mvs4nYeJsrPn5rglgHGtH1o3u/sVoIY+u5WHj3s1ANhMThFH
QBRJb2EuWLuTB9XT7/aVOn3dRqNX9zfCa8E26btz+eILm8zjwU0zmDihKt/DpyewtXiwW+QmfTYa
NDet6dleZfVXyPcR9t3a/xGHGjDDyTdi7LTc5aD85QYeJiGN0MwlJCRhL+ZB2Iqa6wRz29IjyS6N
jA+j2ylwbp6p/HuPRs+WvfAinvJW2wb4kt9QTzpOajdeaonaNQr/QPnDxtrSte29G1CB4njtzJnF
EnC8WsizR087b4AEQoqd4CnP1MYXMKYudzoBge+qRWlWQHXTWSCa2ZMxGg9vtdQCGyuRZaCavfvI
ydIUoAaHu8Ic+PAT86MvMtZ6dv+aGYIw8aO1adF/qFzdrC5xIc5RTp79rSwM79GXioPorM/udQiP
ZMUQP91hStvuez2vZkGZTPuXGW9AHMRZ7CSQ3rUxihM5rhCMLRaaWrw3wf/3m6S1fVo46aKMf4Dx
tZdVyxo7biMgpd4KNgHK9Vd5LsRkJTdKAqrhxb7B3YcPmJysJ0ZoGGqQWStehY76/5Ox3MOvehtN
pi/hUMXvbhs+U6+ybiHW7+EXJXPwXUvIqgINk8Q+CPvayOiL5aUZnvsPKt926X1bYxWG/Xk0roaT
WwtuVOdLVp7eFMB8kF2T4qWdrdmVc4iL6jWWE9GTGVRY0nkyeuPJbMDu83BZJb/O7/dy+gh/tR4/
2yfaLB7m6IYwyaj5cfIcXMEDx0qqWzYuLDCpcqRF/vdAcYMKqejbXaU2qGWOws2x6S8DsiJwCcs4
Cp/ERPyk3xw56JMA2ydQhU9Jij7PcZduZehwxQqAfifM6SrU0FBkjCU0c04IMbKijiNpJenhOliD
NNRbpG7AqpmUTNU4I/qR/k1mVnGwssP7tMQMrSr3adt502yRaAjFI1peTWp3zKxYi5hSJIQa/h7O
4gfPxRcZ8vA0TJJnc5p5iWxBU/S3wZxpNNQlPL7LuD3yoMBpx05NRvrrRfC0sUW11EtEV3xjsfQd
Rl7kT03VZqkUNCEGS8oek3tAHxdDYfbqMjfWTpq9FEt/05uJwEhXTWIugktLT883w0I9NWb41O8k
wqpGTK7fzLiBSFLtrdcFmLywese4ubhlCtJ6MdGBtlRU7YLGQWeMgnaF0lHLE0Su0nQhUix6uerR
g+sCTLNP996d8mhwSjK4ob0FnIs6pJ/5XDLGnsDUexpqJWRqKTU9/+gkXDTomcfS0OzikJCnbDq9
TR2Jp8Q6E3nXQDwSzdOxrzViU+ujBVElUolyYragv/pzJbaTllC0xSWFrqr3pFGLb32sMfxvAjs7
vGtI0Xdw6RCvk01cwe58BY2y//hVgxsr1kssA29p6Ull2cyWTkil9jTnFW+pW1hNcz/FRWS5xpRO
FtTtsjLAHOAjWkF0aobsGh96csP8IxQyohIa5ta7nzXMoTBDPLXdvqnGO9fqrEEdL8alYLNKxpbM
iOhzk/kQgnIVrOwVGnealEIGTk9+jmsZYxZg+1xelPM46lZ7qxECSOfGK05ieQwG6GmZkwIzjp8K
56QI5INIKCF5XPdgQ8KVFSNgtZgnrmT6004s6ZWSZJwysLmPjqjOljtAB9vn+w+fQpNdta4BmqPv
44IlUCJKkvllY52G7/a/JSIhoh6hSaookzKwihJqYWAg8R7wzUV88tdBtElX6AN4gYIyLxBHPZeh
NRTOKMS3NfYGzhGFPxb027gs1kPqiMxXWc75+49ICM+gT13UXhrKVK9sVEo1jhNzx6czz6XS3Z63
q+dU4rLwLVYYcEYBJZgSIAAyOv5Bj+9RYIs3K3h3yTYtefMn3M7C4pwT1Ec27DZ63EAMprMklL0u
uhGVMMguqf0jTQ3g3z3wvrxxrvGZyLWCTRKV3m2r9NqRIfxorVVmoxGl88lQqb6aPnzsLlHl0xdY
HR+dzsll/oa551UZy8btlVJvPyBq5m+/zSQ5L15kTDjx2tBLb6O+KaX4zmi9B/k2eC31eyNffnh2
9xNMdnvz3togbi8Ef8DvFvwLKY4VB9PcUoZ3DU2wRQkCwrgWjuaAir35griIClFzrKbT5OlosTtr
DfBe/Y/4hXfR/VFYeH9yGgoiRIljMMq1UpF65Asqrm2Fv2R5TX1SNDqiONiwKd7HjsoTG4mMQsZU
pLl0/zu06RgGJbDJQ1D/UQugQDHgE9JOHmSInyOMdDulNRnuyJ+9ROOhmsLUaIxs5FYYfUE16WEF
g27mMUOyxju5hWB4mm23H6bxkJAQkpfQ59X95o3GqEojal2oDnWybHVKyf9OUsU0rIIgI8xHWgau
M8KZgpVOWMsIz4lf2ASgyaWihwY4VL6Je2bUlN8KTU09Dtn45KxuElIcDEVfUj1LRHheQGKk0ERP
NAlkKQ8JIOPYYGlSNy58LfKSN8rrIoqJkl85+WoOlItvrYxEP+x2Dg6TGqhtZlN+7lDZrEFMyauu
egSIfU3eACUceTqQQTa9tcE3rqk/SWZYlOORmST1JGQ11Va15ZEoATeJllzHzR19Dq3a1q8Gu2hh
KSycJ4MdSjiFxcla4fyxuh7CM3XRuy846xvMsqAMw2NOXzq4pUifGDWg2nRid3iOJeGJ4S3bcjbR
F024ku0nJw1fT9YjeN00HqHSUYLfv7nJJitg7PsFGth94wZY0l2T3wLep5cDyFvCHFrnWSOAS2aA
6e3VApHQKPoe4suSVOcEFvkkylz93SGZF9GoZB7yTsZ1hP4qtVNrD/VaMM7uDaPGABQGQDQXLuSQ
GtZ45LPiHw75j3nQxyqe2Xcuc1Ywb9KcCd4QDwR7DJBwRA/iNYrk1KuSbFxGqcHG7O0p33Md5nIk
Sui+jsSbqsApNa4Mr5gpMc09rrBGZ18+QxKbAOwKPqvrLT64/DYnGhOkaEfvZASbm97f2r9Y/HiW
7B4Ah6EGE0t1ErwxMd0uzzamJw77YO765qHqbBdzydc1Kt/duOlIxJ6N3GXYw1YkfAS0Ndi+GRe6
02CmOkv2eXaKsjJ1/3zTa+5rCn/sPeG70iq8+ANylIVcjTDgcuOEZgQougieu+o1Hu1/ycxvJSCD
/HlBTBX9FAYbiRFXowmzZ293WBoAFLvFbMNyUZe4hZpIe7YnQLLe720X41B1oPP/HGbMGyDkoOzt
E9KxP8ts7xV7wyh2kstpTdpGdkiunw1nY2bNO3Gnf46t1zOz52+Q5fpYggpZ1YxYzk91oZhACdJi
9D3JJuDYUjd4Bb7MEABthiBroOiUYYwj8hXyizGxcOtgoFV57ViziZ42UH1jeXAVj5XgFFex/THW
yTr2d0NsyH2SD+a8ikqtltI+AgY4Mdgiq0B2VMyh9lwPmrbXFtMePRDMf5+ve6G2m7LH6tHcApax
evETYBS1c2qnyEK8tx8hGW0gFoq5PyK3bkV6o+6tQW1yjYJMMha2+de076Ma3s1oTIZ0xdZ6Uy7x
TZUiMWmA0G4w2bAdhHRqzQ7sJgooH/cfMlvLB0nlMypoF/KdjqH9gA9SDFFG1g5AljivF7WsjfpG
ruqKBKxwVA3Kana+xuUrUDyazYPECLuc7obqiKs8MLGD6YmoQqgizmqcKVNTxJ7SLK/g7FH5nSOx
D2Xa3goqg0XThO72yrdN8xkzkWpmvgOrk5TWRaCtbpFOb1S1FvRcUH2jjYW+sp6/mbNC9ZpjFRBd
mrbd31I7RIe8cxyBaZEHSJWEyqJOqVG6XOHYqZmLSaf+7dc0zO10BuVDXZtD2UMmfyR0z6i2jDEi
pVTnF2uFeoVG+7fIoGcGqFKeDheLVxR09IhHdx/DlHX59bqQIGIFqsLEud/Q4WZfv07lMw35czVi
pHO4H02f4FWTp96LWgcDmCO0j9XHkAl3n4HgzcixebXeVnf4tHfWrt1mIZSrjXbtxJf6ntKUfIf/
ShUBLrRndPIekzaEoNHoXZweQuGYInBb4ZEfo6/bKWFU2yKypllSIzna7n1aAeE0jTKvi8U88bqu
lXsB+fq8cJ0U77KOUpKyNcp+/DCegiEhrrkDaivqgFg3vuzeyZJO80eRCuEG3AQAYrSPmAKusUdj
2duKZUl4LhQYLgW2dP6SW55OZ9yNM6n9DvoHYI7wqmVvyvOl1/zlxiSJNGUWaD99KtJh84F4TFVv
qMBvvj+ENklo7COY3353KFBTHYMa1nBzINGfDr2MBvHxmLbZFTp3+ZKJspLPoMMxGPsYjz2+am3q
hDDDSFteX51OgvPDWW04xxbnJQw8q3q/5DEdA2kNQ36mFOm+PEhl5HKPVX/p4QA6qeWc99S+3NJK
MjKmAE1urm9k4UPCOnYRfR/Ix9mfm0GEVi1tkuPYcJjNDSb3/naFLMSNN220rRdosB7VJ9nVqZaa
hUKC3x2/a5UbCbB6rwZi5VmP09oHC4lYjcjpOSLgsaaFe54or0LH2Pc86Yw3cAMP716ls0B1FVlT
A8zGcaU1RD99D0caowUgUIrfpkhYb5+wQMOkQxUth2TUfqRxqHRUIM3rVnMQLQMfae1TyIrVhrUP
9PPxcTXKYtN+AI6E/7RIL/0nYjwmkhnNiDJpDnW7hE0jqDSsCfjMf+PD/L5rTLZxn8Eb/dgZzeT3
TOZpkokYDsvruafG5Djsacy4VIlnYDV3vjq3zbhcKYR5EtmuWpCP9OTxgRzsSrDYePrHkusxIXmV
xUhJNKqxA9lMv/5V1RNEQS6PwyX2euco7GlpeZbzEjR832tkMv8DLFC3Ywinnod7fqJMKtohx3Hr
1qmGI+QaIu0LBXQFSzYm/7eYayNoovR8qVwPd8IM1iMbgcxc/ZT9wD6SzohAlAKOFZLAFHjOPvBa
TMbd4Sg5W35+RYUY9fr9xZndhne884IA4lIWRv7VMUEGHb9F4H5iB1W2wit9XQ/qqEJHZu8enquw
IjNV5IufIpmUQtkf2B0Mj6w4wdLjiWEa03w9b3zcvWrSPGT0QAvWfqpvOJmXemcpDB8PEboRvedX
dKJ2475i3c03d+ArDnyvU7T5Pbn+K+zixwr9f6MTMpwQN8GbuAlGmrMoLCL+Svp182wzs0CPdTMz
AzZERUi2LFazmQ6KSCAkOzrWMnUj7oF6UfW3Hr48XySelz26zmNOGldURWL/vlM98/qVO/OXizEE
oPlYejN8Tg/PHw/OyyrkP1/Hva5oVi0efJwzqMob50DRtVckY7YyM/mHHm7eisc9zQTxUT/WTEo4
ELOuCZQBrdYFHltzL8DR58Wh4qdNFoX02cynvYvBxHDZnevcz5jqEZAkTKN+n/rhoLnU9MFyRkJg
01Safug8X8Qb5wLCB8I6ykj+pirZI17Daj+C5SDreEQ1n2+GbuRx3KLk8PuD0Rau14mydzf7pRpG
8hRASsH07tWY4zd9UZzjJJvztSHZmnowT2N+anJK8d+pGfCr3EjNVvv01H/9HsBrDYPRtR6CrGKo
7FDex51dDDV98Av65UjTJj+JDHve80Qpm/mPA35ihy4miRQ+6DFV+C2gO51cN3gDnqvui21L9YLt
0wwqtV/Y5GoK+Y4/QUTLxCQ9v5eGK8NmfeWyat1+z3D6wPOK4oxdfnFqb4nEuG6ZSyNQXDiFL6Xg
fPaj5njBm5h1hq9uG0JdkgSvhXmEyk05uf0vo9fO+9NvEsnAsG5qyFvMnTdeSZ553Md0HKHQI6ss
7bbfZY52yAq0oNV+LmI2ItCYBEpEYERD9DIlomrOwOo3JH/Ehqloz6qzqXLhiiUwfnkkkxVgUdr7
UpqR45AyxIEGUuIwqFXLbdeg+GMlzJZYSB4TKT2+iTIZwTdwN/ceGD+82BvQw5S15ABG3qvJVh+6
IIBSKsadVU+mdR+aQaz2QfrXVRhrVNi0+er1mNIWmYMPURoi4TFVwnzpuW+BvL45bJmyEAmApntn
c6LjQ0MHbd9lzonP4yVRHo9XkvSQkysvej0HoPwUlfOdifE2F5UvKGWrfifoDLFXcaB8WxWyvMTO
QZR/ags3mpc711Ozooz0bm1396VBZ8h73HbWD3HivlbfpSUB+32iEFHqDyGlIoVOq6IgHiSySJo0
SinNma6FRvjsUbmFdhXPXRFiSeDc13eMZOnTuYkwBCgOTr6vZPEOxRPgIMfXd5q1NXxAsl5sWSWN
pniaytxYOxmR7kaFRM0f9D2xd2MvCf1O8Cw9J0XaIWh8LISJA2WxJhyvJ+Oz8RA9KYJunZf4Hk+2
9/6jUdrXsQDI85PVsXggClJnvSBZu3G0KyXnKvXCv6DMe54IllwoMyrh0Bz5HOsbQYfoiwydTgNO
zjNdtbW7jqpDkvvHvyjzTy+oXheHgVlqurPxpX/nt6CY+zfJx5Zx97x8AZ/UQU8o6A9pmTL2f6CO
aA/6/OhJDcRvs/kaBryu6jFoxcHMRNMAzy8Fwebb7gMe6vFb0FHHjJm/sKrlu5UPPg/UJfLyj+V/
ZqkktthAyUeta9JQ8bIRl1L0twVI+nkKha801gNCdXMjFUfB059ve1D3779arc2U08orezA6TLJg
ZbLaj12bYEeNVxTDuwGgC1Q/3NNfNusyt0hchbETbfQCwK635NPcLE5tahPqEJcxDckxnoVQ43qz
C6ZXbBCmzp2QeeH4KFoVSgHZRiFgnxovxOIS969WhwYCo5e4WwjdtJ6rezMNW1N0rD77ww5ML05y
C5Xa89iG9ikasiZUMmWWN+3AC2daxMCetl58vgR2DzjhiuOhD6VqjWchI5Wl9VZSExclg9zHkF1/
lcSLgX5fL4UV7HWJePvFNcW8nSEB7EPTV7AQQp6RexIiOyHPOuiM98M0WeI85nYRa7uljUjRDKxv
njlhiLothqz0xqtoJxptuOf+tOUM6q7RNVNOyylJrFTQ+vZKJUPmdZYUgzcIU2UqSP6I2/pMUVqi
acbJPn+y71qwuf+3IGJXYL6SNukOX8xA/vos3emC5nxt3RftIXK5tKQsrvF8AFy/xepGwD3320qC
+fModhYrwxWVTaa3F4GIUJE6WD6rZ66m1xzdnj46ehJYd3F8Q7yuVaB9UvGRg6Bb8kyC0LXWyRRR
iVNYrV0d1qY7nl5OxFBne4R8Q3WqNSm37yPIlFYAsV8Div1UhMAczgFUak4ZNGZZpR6ImvvvxqAQ
AhhOABJLSw09EdOjomqmsYD8vTTAW8YBc3T+5IqddBKXj1P7M3t+FRscB8XDdT2SjvUVLen1cWzf
Nw252AJkW4XXyDUYrx/a70vm6vEeKobBovxS9bwOU+p0dN8Ug0DXPCKycRzRyWArVfzJri34RLZg
huPbcJuLjoxo/AYVgB+QVbXUZpi2Oq982/+X+YqtgXF2SRk/l4JWfKqPgpbpGrVB7jgJuuUP2sDN
EMab+M8K5vzB4rNY+C7VtrxL2Z2iZZIrYXzlS77XaGru/JyDe6Qo5oC/mKOuxqXB057Gi2pzY5MT
mVToeCwstfonOY4AtWxuA9Kbg/RpDGsG8DT8b17OXkYMmdtweEfnkdh1jyV6kT8k9qB5afVBlt45
HqI/qokuUkt2aa3KxcWc9lX0hDDAIeYdgvd53/L2m2R1j1IBhkSXnyIvrzjle7AtjBGr8CIiYLuj
QGPeLf5Vw+/Nv/YJM0R+R8RChDZBbdFNcdtRuhc7NsBBD4wBDRz73Rqp7cuSDBMEW73Ux2EuXnmQ
F+MRyX94vo2BPoDjMr8S88Gkt+abK1iD35rzHBXlH0XyEj9VYuUFKg5ifdcnJZBktYM5itXJwpwk
uqc1VtjONIn5wsV7Ybo+ruO1KDXdAmqYJ2qdN/PK5fgMUVXrj1DEpW+qRRoHwzjgT8irIV0v9ooG
FAy3YC7Wm/9b49QIil7jnNhmUdEDYyB9LVDXyK5sP8NvF1fvY7fNLAw1WEp7f2io9V3Rvz1zLUM5
AlsUtt2y4D1tj42M8AmvoRqcQDtD737TB7u/+kDGV+QrTrPyLBDVvp0JC0T8qPloGOYZAHderJ9G
XhbodufuTXbjsgWldlzd4xQ3IIuuBGScty1r2Z7nNaBLFVcl4MLPnvlRYWqHqb5hr2KFblDwsKYW
glrzWns9H7t6StgZBJqB/iSLG/xVvfJnbRsiVUpLTZIwliI0kUed8+OCycMPdbDTEp3r+3tyUupy
MOR/DWOV+43fisz+ReqrMwWRvKRD6wTPsL4pPwnE/lCBO9SHYLnd0C793c4o8KsVd9mU550WjTYL
367EVgNPZwqsz/NSvgiMNXAhV+Vx/irvrby7KCgIsID93G5q2BBN+aJi3Yvr7BNznAUAsdqcIOxE
2+2YW7OIrdhzo+upvLvnMBBtHXgEQZoX+jhCJ7JrHnC/n5FFCGAlfHcdBGvYtygsFn0wvPCr0Cyw
NhJyYXWATo8wEZATqtj1VYrXIse2RDd0XKWakpwmlYpgpU1hq1AdWPOcmcyipB8nxUduuNNdDFZP
P8fuo0UbgbmiYuc76IkDpaYLYbD6GHo83FOWpnxtV6Hl6TBJ+4IOIhnKZ1zU2LeZIkUplg9T9ge0
brA+DPNbfJK5u8kiMRPaZVpfRv7tysfuq1Eu3VZ9DfQgFXFGrdRHbAfKS8BweCKvo1E/OWN9KMk+
oe7+fg6/2DvwwhkaQTa3kWUoF4oxOSsCYju3zzAebHQ6NcgWRuJju2588d+0ori2+IRNd+Xwc8ed
9/grG88ZIacsMe3XE5izHqMH5QmEi2jVk2zYp7sSx0WvuOmpQ0bpimsLcnh/eMgm0qM5seXt19oJ
1jXzVJFZrWbyRsVPrS9PFrlJ0Tdt0d/29EQGZgHP5eUtm4+EzwdreaJH64Sx/Oebiv3Mkk+urvhw
uq6jZZKtvAX7WpCNBavpHffhV6jP3vyhfRNjzxFdiHSy9kdIN8qFH7MSGj1nAZ2H/bGjsi6lt56w
tmnImNaIYJp3OZyrKFVSUJx187+vHaZUpIUoctgn6H5uQava/sApITBLBnPo9kZPvnHNk/HyjrfN
5mHEKXsK6Gdx1dhqZOxsIHgtDcLvbIRLRrWZVSV3cVRz2MIR6XB+7jRpLFYYqgrSc6ggwld8cmAJ
ecMJzZWkLcqpR9SjkjF86az0rq/RuqXiNsMbG5cYS28aqBBcWosQuI7JntAr/N7q/vucfc3dYneS
8X3Un5fGJ2+M9PiU7wxh4misEUG0b0yTm3NIIt2NdYu/f7FZOrRX2q1IDz0732UN902WYxhSB4Wv
OBp9v8RJQh+SGB1/0SdB+lEi9BDmViHNDldeus5oe2wQuxXAH1vxmHmGgVaBH30mewaBdYknAmOO
2KyzI0tkZbOsm1tI/sRQorWnaSG36g03ELhMM0tziEjjInVbn0mURFr6a6xGkKEmp9N6WD9u4gJh
yxujOm/DjnYLHBJ3dqsJVPFRlnnfvGUJlrT/NrDUwU2FfDl/mABUGZ4h8bQjGueCF1WZPaD2I1ri
nWV7jo2yYMRE07GIkQctGlhcVmUlXvIvF80rkrndK4HnyHd6xsyZvc/s8LLOS0a8hsNf8NZFimPb
OX5e+bF1FK5Ha8wrmlzM+KFH5mFxS2I+WFLKfpUYOKXWqNlankb7rCwbB3ZVK7+LRBS/M64b8Lxi
HeVQuEBrCKhITS0eyMhBEHB3+ZvL1e55OOBWFI4gtzlBY3WC/JoPQGVUa8E0+ynUmo10htnD93da
9uM7AsVHqZ9LbH3TFlmCbtkBfEiQN/3SP+XYYCwAXPOdCuQuCYzC9UWQ8k/j761RWXfYsHoI0Bpj
4kVKQYlOMpkgPxXa7N2OnVfAU6y0v4+C9IW70wO2Rcpw6SCf6pfLZDJQ2VV8U/bm0/sVvVXgFRyu
ol3CIOgggfP38M3xJin+Uja273/qGOM7tuMsy2u3u8lhnbR5yTc4A2bSjAFIymceitI4aoDu1nOQ
L6gfd7OqaJwslT/rV5pV4r2l86BEI8Y+EiPfTBQqnKeyEb2HJaBZaWTYTcFjTHbkfhfkqySfRNnW
qWejfFoO1jyKm6fz5twFCN9F+rw4yRqjcj85gdpj84m9AmFU0sMqHHN8FOm6ymmLUGO5QBVEbrlS
7ghQfDMVvQRgYkBGxn1XGSSewcvZS9ITG29YPwtqrKzRBNtehNvSWOGeLjHOyiTEFiIt7+Vv0X4y
cL/tPqnll0Zc9/1YJXICR4H3JMCx3m8p4RqsLHPnPKJ0S1L4zC3vhkcJUD9ngGP1AWlYPXIbrS1i
AJtEB5m76soUkgaiyM6M7OlMcnt1AsNIBxr2b1n7Ktyav2rr/nZyQWeG/qwyqpm+UIi68X+8tadP
Jr0OvsSyV093azIbOThXi1nF0Z3uqPJapXFlELxNFK37lSROCmaIiqJ0dUXx9wMnCpAbTwMM4hAA
gdQeEI+loS0m+4m4CODIBsYygtVa0uII976czVRPD9+TCHMl+jB4GG+Hw4VaytzhqaBNb9JD+Nwl
V9qhBf6exaBQNTtjVJAC3VCblUZhrpYr4k9HOHSLkgwIgpLqqcB1Dkqj+FvinLxaHrafCRcikfk0
a39vnODkAfTjExllrPd7mMeNwGzyvXzBWcP/IcejcmAjs4GbSj2P4ZVZAWToMLrE3w7GhFSpmLVA
ztOElgREqV6V8Z1hCC22JOzxM8gU84DhwH1/ErHyF0j11xE6u28sr9QprhPt8io+vAc26fnW2zOc
UPjZ43Nad0qYO8TSvwcoYZpj9JM81ugqgyP8rRqZIuAuTuATbU/2dM97NsRU8Bl1xnaOag4FkuNe
lmLtu32sDEheW8UrbE21Lj/rpVmnBGOYcwie7a1GqexV7UlURrSfATk4OpDWz59u4WuKdxvmBQao
zmDDt0tn3+S4PEY4ZpJhMOCazluXrtvI6MKGd1O2s/hG5oxyD604JuC+c5Ejmsw+DO0eipknghe5
AsLvsz9jxqG/ep2XoT4gQr8tee2Ffdg/0CRO3qRDB3jFnp1vYv5N1ZebtzryEZ8Y2L5RZYxHNJyz
UO+5HUgIIkWxWLCUH8Et0FI7g8fqjICc2oF4CIvOT8QQ26TjPFSb2L+pOS7+kLrQKRRGEjXg757i
OeRl1PToCU+XoXRBzSLR2VUGTYs1zvf17D9L4p6tyo4TKdWlQiVPaIopW0A68KKq7XiWiDK00sYn
PmZVpcmG9HM/JRqfgvWuJlcjzkwr8nROH7049wQRjZlsCDY16wWYCNpfJKJkHKsSD0byoiORzyh+
+iLUYwakLqTQ+xyzsvFRMCDUvdwsav1gT58TlZ3AyR5QXaMbzRXlD0XJSAxuX7+QUhL15fYNWfn4
+KzyGF5+w1UqesSeNBOSO8a87shucroDDbgXPvjuaL7MaSvUyYwR2Q+NPmoXTYXGggca4J/2t+n9
ynHjeT4dw6YKNmxqiUuDz0FGacFEH+VVpRCC7sjxCuDRRWFZiAB6MryzuPqHqv9F+jUNBRVZHZ7b
w3QZTloF5q29TVrYbAL6oOSIZqglZZaEKN76w3RY9U9N4AAA5ID2BzZEQ1FCkbxkT2JSueqLCPXZ
YecfiaUew+aH7RUZNj9yc4ymX73+vKCxhsGoqfBCUgAhstL+0q6vhYS8+vgT08YnoLjcKKI3tnJJ
QJ3ow3ylX7Ss3k09wWD3rB+hZDncEUwiM47pXRPsZzxRkxNVNiTMxil6kXdgAqLnSP5tmpPtnV13
8Za6PHmWf3yd2fy96wrWgLk7txgNZRLkwBPtPwmkuoXn8VkkTT+mA2eVir+JGrdt6xaDCf/cczJU
NkmME7sCqlEG6RLB9329V8KV5Wvwf0s9RxJxB438s+hf5Nz2kod9CdiGBIrwHe9SIskuCgrREPG0
TcdH//7YC3CIze7rclvLOC7RAbgySOw/7Iw1hrD/CdEh9t70cdzohrtcqfJCEKfH47wY58q2Va4k
paOrYBb9McgQ/Ay1ukHQvOGSMGOXB94WywJyjy9QMunsnYIEGKl9oe8SWAAd4gQN5owvA1KlTz+T
ofF5szmkSg30xKgj6ALzPk8+UojyBTxo+9XwBeCZIulUHbVdguuZZV8M+8hnAzJdr8NdBgX+k7k2
mkpHwBaFp8gpzN3Z7axl9QSaK/RybRcsELr2324zfCCPuVWb3cLjs8LRR51hsy4e0+dHWO7HG+g8
MrpIv7te5sbwP59wjEZRwFn74oL94jOtmurm565x+V32kQBLHzvBL/6eu8qCGToU5AROQlR9HGyD
iMOn3+meT/CbdAyUKzQGmxFV8w1GdAffSbuR43sfxUVZoSkm6udpDwTZ1nayylNP/kLNl2OTAPCz
w8Cjfm6+P8Y2mUHZqO8ZPBl+ph1xxv1g9NqaJvP1xySjx6FYc4PaFMcRjclHedKRMadNOAaKxaSS
K6kSU14quaoVA1/lc2BFJagDF2Nv5dGu65bUxcJyHMLkguA88uyktxRyomECGkaSjXQw+7FSLcYK
twfS7GTIpZQUiHQnUc9Kagab4pT6/ldhuqaaKbE11mfFhgONbVkeoeQm4xnc+6R6Fe+L0pbEWgeE
C2iL6DjxnrkwVgEOZox2P/XKDAGHOY5161VP67ihPQgoQ4xUovt+3dPTWnrSnh0uXybSVSYnTihb
HNyZGAyonhR16/hrfYkiRkxst4aRo5TbOQpX/JZxkcmouJo3mQKWQEBaZvetsPWtV0cbjEGZvqwR
YhYB1Jxa6jFhKGRoG7cJudxYwrECYfcRLlE8a2Q3OqwZ9BxzN2NquSVf+0etKjjGSfqV9yCyV1t7
LDMwe6ST7cw+IHyZvfRdbTlAC6QA59rb5nhOWHCJSO+tD//kVnf/peXRWGP7F6xDHYEO1qGOI9CP
LWnGIxbzmKuQHim5SBSQAtOmmmthM70+xoMSVZ7Je+XGwgfp2i1uhqo/XyEpOR7BGiVjTGHoJORt
F4RzeOaRfrFmZufqnj5b/DEohiVScGqAhpaZi/l/daA0bIb3IHLFCMlMDvFztHS2Ms26ZSwhkRa6
T+057OBJsF8S8x39xNFr3kLIRclSZTrTdumJruqy8l06Rnj/WRYD3PLAVh9Zg3XElH4LpvlRbkTw
nv7aPJ1gUr4g2+zQO+eOYA8nutJne90HliDqXzDvSmzr2+1o6dMFwBlQCSlu4n4c0ax7mlbiceHR
HFRDwagRLmKH0mwkTampQzkWMJ3H1sxep6v29LI1/0P4//yZZE3Dc2XMsUp4yCdbUqttT56SDSl8
G6CgNeuaPXpiYvfVeeFyVlgutuSZTeibhPXGug5zgM0vM1K9qMCOWezJ1P3ACoSSomD82jXani6+
dSc5VdZOJr7Mgmn4xg3Ua6zQDS0VbJ88ItyMnjeyo9cBy2dfM/3q5C0aBGR+9qstKbQHC25T2DWZ
2LOnA+NWDjpGfxdftZEIeeMSwjDnJrcWtmMTrrdVB2VXH33oPrIfKK+zJxas4/38ItM++heKFes6
ddNwX1kwFF2rI1CM6/yuiXjgm67NKL7x+wNGp0HEHW0UrDq7ZT8Vt8JO2w3vjTDNUUdHlcsEwqSh
PC9wkZWN8BZgZEufvLzLKRQlpHSnfraRyRG/vG3LMhGkrYAjKWKv3Vlok9MRsOG5um96dKOIzWsS
OgY7ZmvdDDJ4BqHMhhr77UO1FRAUwQzgvtQf5SAo0U37xM9dnwijGeKZIiYNDRdz55aFEI7++3vF
ZG67TCCpZ8tJuyFZLE4mvNBo2qQMOXkh40g7kc4ShgrrkpQ9NcHFAh/R39BdQZrXUi44oymNM07E
P1GgXg+6HwKTCd59Y6qJIxhlU2r3rgD6u2uXtVllsFOpBiO4pgZ/ZIP/I2+88+fiiaX5RQ028cva
WLweobf+NhXT+BPqNaF81FGL8AyB2i0wer5JDJhYRiYFFRKU+wSTAjoMx2P6caxLie/OTupWWRK0
qpilWPy3GbN0lCDMc3kLW4NHSS48IdEazfQ9buM6pDPjb+Ju7w7Fy+WLRDkfQWaQHfvm6h/l3CUZ
Rq2N6RPTo0pmNQFzkWgeDZUPWFLtrW49XnkHa2eDY6obf/kMrxP1wM9OV6hgKbboDUFOSZsdmUVc
wwzRqy3OSS2qiamY3SpbuEt/WHZU8av85C9X6VHgicVkFartFh2OCRXYU+HAMpG3Yvuo6v3Klzgs
n2tYTEydxdEFJgMveNSBhPwzdPAW1mLRZYf0cnAWt8X6hfidNlN6UO9IgcXRmp9Qc5uc2WLoeT54
BpjpnYywlaFGOXdDkGQc5SyUSoePmwsl7gHQh8aJ5FBN7lUj+w+D5h62yJ2QKOf8iH4Kc1pFUNyH
j6gzvKacB5v18AsJMKyE+azB1IsXeNyYbBRWIfdMMjzobRQqlmsoyDcr+Xj3SElMKu8Tu9sG0kxg
AV/BeW8fAiQuDXsa8mL5YQt+Nj0goRj9ByeJhdRLsojOXfxfkN42F1kW0iqlKm1Kpq54St52ZQY9
mA/iXD2vSlUtXAKJmliSUuWty3l3/o7wLworKuvaLtakoMMvnMAWr5bcKnCPDUb58nkkOfAAfoLR
6Edrf42LFvwepU+o7VGa32EnX8bzWkgnMfYn8eY1W/kYALXUBXkN4TybQlpfFp9hNrm9QjJOXs01
cZfGigOyWPtk7NZMZ9DuOY8xmL/gDLDgTPVgsWJLgOXEdXItPjIRSX/Jqxxw3OwOAIP2LQXV0MUI
e7h/1Slbtd91WzsAgCCzPPjA9xf8mlwJHZx7hEHvN/9fPNHdL8fz+yc0ruRzqDlx2OgMVsjxNqmE
L81m+KsUmdBrIOaqexSSJK8mydWdYpfgv93HG+YGXStoQsxkpm7u1kTNGZiF3nwuNLxh0j77k9o0
OUK56Ro/skRRV230Q+azPkyW/VoLTIvkk3re0GIVOJGq21kExOJk1FTQJ5WUr3nBUZsZutg2WNNC
hownYiTcA3zF8q1rkdDgwN5gzE2b5IpyLLk94rLdnvSuCPfZh+VkWFeasItXXM8Z6lykNmczu0U0
km/beeuwDh1WZMszsEh/AQY34vODA0FU856yYl+D8Tr4OW82ztwmJqlcrKzuyYPK5CjJrw18HCvN
HzCW/0cQTFqGYEKMb08L5F5vgkurUOT+c0yis+c9RpcSFqYCN3bTiyK0oszjXqtew833yAfssrZ8
ICNO8L/VawSIUX3ifstojgy2vzG/fuunAgSa8+BRw6LyQufPgj4Wathpxi05olUTAzJvsW3AwEcD
e7yFxKWBtum8ji07DrOWq02i37+emdGbzb4qmdyX6TIWzKnmQl7BgJZcKhob7MtF0CJUBXGQX6v0
tCBGuXtbzcKN6Fche1YfgVVDb7HOR6oGSvHbI3HvETEbm0eySSOIIfcriIFG9YXRvEiCdYKHJNT3
p93/h1ion3ZSezbboNypsjMapHLxZTHRxUoEIzrLdvfOtEuohfXzkYXz2hJSmF+LLdkOQOMf9OLq
PthH4dH+85xX0zPRpBJ+jrduLuLXWMgIXBKWqOCiPlt7TQw3LIcmqfykR67v4G9miSYQMB7NURrg
YWmPKRWniMgGqsQaxokxs0WotngmHO3mryjIHVCknis6gBjffBbESFawVKVRMucc2+UCKW5IflfO
r/2fOc358G1r0/Z8H3J/pnCf19mr1cRy/LQEaoQt0k+nfiGkaZUZS5kpGzM/ENaK2hx1LkDqH40R
Y2Sf7cvcYLc12yyzIS3dXgkv1MjSY1GTCEPiA/g1JNUnnx7mBxqCuTmH+ITQlLnGMgDNs/4glEvR
Snu0HZHgRgKayyxVXWMqe5hyDRgzEjDHAty/4ZpICqVZ5ri/BLwjn5xrEKXu53/2TnyBQfp0LQTX
L4ZavApQ0vhfeilAOgaWtAAPzTDwbKqZi4ARaScYqHlHIrpC3M3IcyG6KXO9m1QONLzAwU+Vc2N9
MCvmReSKfc7nIAh9koa0DCCX9XvhwYg+P7/A/MqVaepGDev918ZXgjeOTnvsCg9O+4yUGGyfHVh7
W/0v3anKsa8M/XD8w8RExi1BjH1rOb3fwdEBMEo/HeSaadsiEb4Zwp19c1TEnrWAaAo9+/WySP4b
br8GILbsjyCf3CXYId5TZ7r3bw9PULbFEKOZZmh7lbUgIavbPDWYqN87XjarL3+PODFmGqBBgmWD
BYJutosrsEPuaDc7ThI3WaUr+jhzJK47ntc3iBAfWpjMsH/IjB0vINUX8UC3WORvaH4oFPk7vshr
gcWEW/s+bvANn2Wwa/LAeQdzN70KeiQeePddL8crSKXKLiOF4h4VFS0PqB8C1PpbkO8syFSC3QcK
/Kv1BI/0euWI+JaoInbGZVllZLgQuhXLMRsOglwHPElAmherwd8vzu02IDVdPrRfh+/BlmH+HLz8
yAqnJ4tDP+jYkliaitOfOli0d0WZsReiUAhZZj26Gg72NGfqTUyhQ2wypSMUlaSCka9Ddp8oJ9CA
p7dKJ4PH2amDRHfwxdE4Kfari+ObIyd74DJOO6XTogCmZNYiNtzJ483WkDJ2/P0tXHLmgKeVvBgk
m8cs5Zwk9IuxpuqiLhlQVyGcistmHmGjlbvyaXgZTV+IuiqJ8EBgNobHs23aeOPzTjjIZRLkL6Ip
B//nch+dbarJ6KM3jk0v8vaBXvkaozXRVLBFaZMr5slJHRpy7pZlPDj8VprCbsk2mYIggDVxK/gR
wvshYY7K+oqgCfeTST3sDqgxIsTryMIEMkYekEiONW/seTpH0STvvhfBMUvVpYPtxpEFAefFFIDq
qS/ui3TaJoasWJkP6U0dQji5PZhInGvVD/0bkKUBLfPDvfziqvDp2z/vqJ060KY6P9IoyOfGs44w
JcD3vh1jwVIfx4TGbrw9H5+CUqliWrHZSffi+5/uXmlRGtGhheo7x6UldmteJNX54w3w5u9QCL86
qaGqrT9Clx5idUVBj5FjbvBctKv+r+yx5nfocArQz90484cdTCk2hfPJQiDaMI6gmwdifBHUJ9Nh
SqcH7LnRzDioK8IetcQanv4WI7ONcQVEpH/wKVqbLV0d0/MGvoovC1FBq4ZSdUg3yFvOLaR4XbdA
DK/tLgyP1MbBLX8vNSLfWHvIZH+ASrUogvSVOqu+ZSSLKbgjVMu8G/KjLySIknmGLfs7GDGnO1rh
6v+mAG1EBKIQbXWNp+92q6vKjo0xjuSmPIxzSp6jvU30IHHInt1J2Lue9bkKlhPFSpRDUlRpUpzt
fmXqKhV8O7lEK6FbHpRmwocJFKf6U3SHwGsvy++fVenDWYn3MLoHMMchv8x16x7vb7+lTwLsxT22
Ye0gnOTVDYgiEhmVLv9fhrHK+e4LHaQaub7sZFfW2lX6LpBYh8TeovwX27op1PuKDmLCa1e0PRUk
KXyDwGCNA6ZQvK41NK0mxmYlKvJ5uW9O4BT2FosnL4D7LnpOL0/a5geFl9r+yZH854KpuSAdqFM5
d0Gs576UtXrrr11iZXKH2O69NWBFvkFg1Itbj8XxPCNFpma3JuLamNKIgXvr8YolUD7UdMl1pCDr
Yk+ItqEaLu4iS2MAWPCB3j0qtcMbvQhAlQVMdqX+TmUrSMXLEtlKljKgaJPZ+igiK4ybHIdy+i3u
fYAL9q+nrstvM+pjisI9H9NrNfV2WHnuWSynKZkpxDW8oOGCA6gznhS6r3xJwESjoqU9V54xh17C
FxX8zCwsMNtldgkQMnEJ0xobfKF9vMvnjwDavji9AzrHAHwqIn66SrpsjmdoV0DLk8LCfTA/kLUN
7BpjYETAYhyrO0FMhqwLIFRYV2t7bxhuoAuFkdyt2cb4EH7/3hXlxtIqSVWfsyi1kla4GUNUR3VN
/jQhD6YBHpq0RusAAvT2Ja71uRmsEvJ19/UPi4PacEILwumDyqDkmfJ1DzanpJ8685gmnktvoDXP
j9XVwFUE9PH5tdOeoAvGa3v0vKyJ5kB3nh03s/akdD/MMYyh37G0CG7qiKuVr3ZQtdpLsFXUeTFj
z4w1S6cEx4J9mrYzEmWF4/ujs80sc7AlDXfh/5qlqtf+4uziCU/0+A6GNUrvcOfxUbv0MumztPa3
ACqbXRjCdCqUyHQ0dYCAt1F5UrR6GCVr+lRKVGZwqVH8X3eVKU8QNwqvZ/kKRvDe5ktoaK1HjY1f
Vgo+Q4789yZSGRK6SXrHS3c17nqWOP4pwjNA/BdT5yUWa6YoZ0cZ4z47++9WYShdFqhlvzlk/IYX
r+mgdtDjP+cAHqQAiAO6Z7URGfymOjnJ+LCMVXa+ZPdDt2DU6qRuKefDkXeGLoYstp56z8JWk9T2
yS9kEG4bOBOUvv3NMI1gH8mWgIjFzejhIJmy8kRAUNfRE6DY3vKSEgPhRbDEh5P3RxIZ62BPlqmv
5hJnFfUQtLmn/2MaFSW+3mvG9ErPWwguBKtLyPRU6NfrZ+mWkXRnZL0GugkZ7TrQHRIHlZWMDadV
FQy4j5tYFJHGZTPttEMU+PTrYUepyJxBhi008AqQs0hHrsr5xWEq9ZLC3dzycTR1sSJV1ofwvfNb
JljTsxrn8r+vzSjGkmAyGAtO3Uf+SxRjVT46EDtGcJgcBPqqS2yE+WVPEgKrUyDOVrlx4gf3XYlA
HTCDWaUErN446vXHchOfZJiJwpKjyit2LCW3At2aovsqA05zmmLRm367H+sDg6gr/T72hFde9ldI
tBS0GM+pTde/GLJ+VjW9tSlnKLArmYUwBNS/DrFQYmYQM7wGIQKBelxkQySCUygLzQEBytn+M3ps
If2AYK0tgbyrOk8AHWo/8Zw5og5n8tjb/iCkl4pmn4sAC7JIaDh4R+hICzV5Uy3A57zpRGUq3uYQ
XxEccIPDZDear2EBPAei/QfXJ7mrr2MOevwL+iGtNhiAkrZxY5Eu1s/UVLMmngAd9fVNQZ8M/QZ5
wZc70n7AJ0sIrAB2dzShnQ0kYuOq8Nx9qRmIJxzcLCW20ZsqYeenPWKUuUr1zs7NppQbCGEldLat
5kKYukiw9cpnHBaOKKFiarAmxiIwvUt0H8809Ot//laG+QF/0hnn4tWgnXrpJUNmr8XgO1164XzB
kDhg+Q8ySIxwW2MPQZhimHZPkzud1lvo3+UY/11cNh1gmBmAKD5ACqfUnhJUDrDThb8xI2u2CI9X
fRiGSTUDSkh18vqWrdSYtj9KH9a/P0jfR8Am98g1pAXDEC82GaqQKo11VkvLlzDfkcH6aZOYXQGl
j0V05kg2UJmFJ28sPd7ft1TIXF3mv2exF+ACJFSfaMgxYWLDXCUePQ4N84L7Yf+pxR7VjhYqrG0K
ly9JgFu2On5mi6flhO9PHSSW+fSPUcT+ciUorYDK2fAyD81dx5tWy6cEGlcdNArgAWmvk3ecU1iY
NaZndsq8e/SuH+K24GrLTagb1H2A1p/Wg01OHvShyDmwT1+Ib9Kjm0OGuhuYCYpwhlRlcozP3IsJ
Y0Gqr9pctL03xa2NNvqw0H2s0iycIcQB21Lrf7Z+Q/DrRnIwpBRr9I1CSZWHKOwwrLf5zrnTW8Xe
UpC5OZtD5FxqMVh9OxPHlj6M+PViWTvbu9pr+lnj1UbAu011O8NkipKSxIczsiCWJ5X49PtfbnfT
OaDz9m5VFRTIN6cirW9X7UAQuppcyKvEJE1apx7+ZS7oXObtiCMsCLJRd2UsPKsb1G9BeMvmMsej
qk3cD0GI9BQphVjceG5yd6QCqmJxTUPoRce2xPqitvzDw8+IGLLaIulpgXoFkuB6t3yTLR61Ly7t
3PydJr9p2jJ3xwMiVmjmXT1QB0aShI0mFhnuYshrv/VQgPPRoCzuuRVb1dCMAIJai92UyBA/0N71
HLdO8SMBrsOgWWGp0ZZma+J+Gw8ZL1mtEVULOcY18ZqtKsSFpSRtQbMnIbgVJX/Ldmg4WGseRUE+
+VHIcV6N105DrqKK12yhAXu5GDnJzY1q2WSPb/xWAIrzC795Z+tBlar2Z0Kb4FBbzaqA7t7mw0bN
nHLoK5cSpi6EM5jv92aLZbtUsA96EaL9NVjPnnw1URgbMVCfGUHsl1kDMpL5EfbvFAKpLXTegjO4
cOoamXZYKWKf1n1+9kAffDaFzF1KaDfMRJWF+bezjZpDZ+szShkULP28Cl5oc28Gwd7vRjKJ0jeX
NbotdhJTIJIcWXthwezfuACRzeQrxKIiZuTWa/Fhn+vP+BUJiqOt0VPgQwjHhf+pkCjI6GfJXi2I
IzuALlj93z10RGwtOIsE6tpnSGQljG6cFbpTr+pdwHQNrxzB4TT427b3NJeYsrFIHe3+mgmj4CCd
WrqO4UTzBkNWCyKr+IZzq8BO+i1OH8xbbbzaH/87EJvoMWckZKSRU6S1ZFGYQKROyOIno01OitOA
POZHOcHuXWxhpqapgrfFiJOXGw+BQYTrCi+UrSqIZxbBq2CDpF23Tr79ivmKtoJ9cfx1NJz1WFn8
L/Fvg6FjKblsDl/dYCN83SxISVyqdF68uCa4CCalAJk4qR1FdtiBsZIHRFzfING3PAId+/lrzimU
Ns9zNdwCvjWjLhOM2Rb0GPNZAqIYGUIi0k3KkCAxQm7k994pHPU1QpLd9DnLSrHvQNAWykyqGDLS
cHexrB6wcPAeJoldEiSdeRsziX1jsK7icDDwzhbqYqmhWPEEa4yCJfoZNWxg4GZ1AVgv4aQfWe4R
R9KsxlCJg8PZoY9kA1lOXr+4b6hFQ41fzi8wfwBkdOcihRR6rNStX211wwzwyfRjHm3Oj1+SAnr4
fM53dVvXhTHKv2QgwIePxMXoUJ/UA4nf16cE1wWEV6hM/Ngk2ZdcO/iOZw3djTQVAC8wNgaPpVXO
iLOBbG+UJ8VhLDA0vxW4+0XQNVrp7/uL9zmMfyfrinLJigm+DehcWdyHbyclO96kVSfNExgarKkE
tPhXnwTkxnVX1sMM9TUiHPN4bZwhP3WxdywLAmUEwFzIWgc1bN8vFkJIvgdHIBLaijdJ7whitJqK
aRpVrAlrcuvMA7dl6dhkwlWPb3s5TCloCW/Q+WL17S50HBActEffwlS1Jhc4w06sA60b67MUkXRO
WATX3NXJY1LDz81Ro9lL2Sq+nBRLywIy9Ci+p10nbm03YggOPUznUwQCsWN5l1eZSn62KL0N8Ooz
xTduVAnNKX2uFbUxJzC/gKe+z3nz9rYJZEVDamhfUJ4LWpfMOZBftXiFIfYZ254Pzf2QRoxb/r7O
5Xgg95Eynjglg+Nlb/D8jbSt5NLqfa9N8L7pPXe4gyfk5tqg4cAsVzeO9hABYhDjm6uZPrsgQDI9
wqBmMkEv8wtAX4VCIat6n2XZhVQHGhqGlCuFnNT7ZIH3mTF8nHbp28/C0iFyRnGaRwJ1OU+nHTti
/DEElgjETA+Ge0V5MpHeQnZm7ZxTyyLo61h2xcmFyHLkonC5m5jQ01Yn6Un5Y6ElfSIWrAEwr0/w
L9bTN/8S8m81+u++En+vR9mCqwEW+qkk6DUTy1OTF3Mn7MRfZh5R+5gHc+/qcbWEmR9uX8uXJdvS
ELJNMe8PtlkSAFMDGkI1wSNbhaXXW9J1lSXf3ld6BsdKLllymp9H/h4pQAvjyejzqi+4M6v2dIuJ
Bm0AEQ4ZsRpmTB78cC2PxyKg/wJvxiQpniCEEy1edO6Ju4oSsiZif+Bh4pefcX5tecG8yc0yAzoE
vxpkIjXz4WJtz4zod7sR1MbFdfM+VFzGtXgGEwL+ZaWq9gwJFJO4N4eEMMdf7LJOsbeHLReqTCR9
0AwSaxZmBzMciDig+vL2Eq6v28/LkhirrZzsWLkHd776etJtj7c+5GRgi40OET0Op5Zj1ZcDImdA
JJCA0pZzwdc8cFNqC7xCEeH+XEa9ePsoh8+b52CWclVQe67W2EeOv30IZTnKZ3NYmqGUAYUz9kHG
K2urnge01Qx8EeK0TBm2/Nb5Er6NNMut2j/LoCaBx3Q8af2pz02CtU5rzH/KLQX1AZDbYUdr/+cu
v+JyfBlQg0dhTld3vrpCs6YQALzvEIwrKFCy1lbuZ7Ude5x3Gm+3ALUF9g9bba9tVfXO4WEABQl9
r9b9hRyTy+IZWiLGc1F8m1TUIerNGXA3naQyd45qF9czU0WM84Y9uwrsW7bHAxQsU63a5xVcATO0
M2+anxckGQHQKMvwFssIsSUm1ahPezg+a2J53zuHZivS8qGFZYXFUJUD10F7pL9SmUnaFQWqh3iL
jJQ3fgsEEKXuhMs+M93FC/8Me+gWo8QO6ncGsFFv1as0ulIuz4W1a6GL3FsQPdWGeL4A9vi1Bfwr
G47OHXqcDs8RY6rkt3q7VobkPSuhCplD0L7+ZUzBfJ7OwIWUmS77+Nu4QLnrU66zxTocM5uK2CPc
FW1YP2CnPmakHmT4kYTMQTIYJTdE9LaHsmjwae20ze2QhThhkVfZWG9nk68yjCNQrMs8B21FF3VU
n8PgyX6HaK1rGsLXi6m/42JGgOi2z25OKgt3plxu2vVdt439lo1v6ng0oKqpYZT3l6efNAETlNV9
zOReOO3SiLBxUlHz3+5uqa1V+NU09FPHFIl/pbtCNio3CzwAN+pBxWp6h2Fxs/KG6+gYFopcTWVx
lDtR2LjpRTyLuVd1e04UvueZeuyIHq2ztPcgM1XB6v8DVS8R4uGZJMXKf2vq9j4bdug42UdLperf
xoj7Hqx5tfwGt+shUtI60f8Da6c9I2rGvaEoph2vbNAmQ7DmfGAjXqNpII/OGw2ggvE+T6uaNfZe
5o6bpQDvQAeJ2l408JDxwf96ozQV50fwi5SATUECA8ow2DrftxgYrfwstewV5sx7MT0AP7+jYW4G
MeDdWz8qCT5CxSlKnwkaeI3qpvw+8evN7BUAFCU2R0sZDHq8ef+X+hjov03+0hmULuj/aUtdQrYF
jXHVk3QmiLdSjdAL7W6eSoJoxMf6ULrj5BOVnM00P9e+zKAufMvtQ+9kYq0eDV+1C5DZwaU5BTEh
/GSPsmwvE93sYDsIVXW36ohiTQNFXUtf6h3L9ZOafdk4TzPpb9hbOEktG1oGQG3n65BxTg5Zh/lB
+eaRiIat6Un+uVtOQ6IcwT1IaOS6nhIY2EhpLPqvZCDdCh7hd5MLU3kcY58DZBsnzGsQeCPfWFl5
wO6Mn3AgDPmWzJoh6uWOjrUW5DnnFOeAeHrvbqKnzKVM7nGCvpxkGGzWrcH+UilsYQ8ZeFUvzLk0
XMbGo1oKQYMJV0i1RQh+Yr6T8MMH+7hSzsPgvwPxSmVOkvuGZ3BfjLx48rCeAgZySSPrPi77ojNI
3FCq5b+9DY0gqfvWTYvENYtE07AfR0MlokvWzFqOm4iHIuT3wTTTPaTQktaOSSDB/kOqdyEnakV+
sgt3l7kHRdlnuVe3R5Uf/1wqSxurgJ7V4RHg9jU4AsCSi1gxfaUFB+AZ1EN6jM6UaDwfY4GDtjr9
paPn8GPpSZ/i8NWkJ/wDR37TIJQB9/7M0wgy4ZlOYDJtKiC2Wsn1U3vEC3X6ZKF1wH6GBVXk0oOt
2SKoxK0JOUn5cD6UDugFYV73mWDwNofeIjdBLbVA5JXMR7Z6kEJ51d59Rxbjys782IyQvaIdnm1E
aaq3zKNazYRjYL2xcQte4spVdOmo8lAq9u4n2QF+PUm22wFXIB5kwLguqBkFA6boilQ0mxBDHZyf
Rx9YZTYLG7pZUhbjp32CKx1P5dEPGRsFtJ/1poWIpjoemWBoXm10W6Hkn6f8XGW38qgt7oGjJfVs
HhoOB9joGVHPeWNIclfuUWCIV1Dq8CPhnINIkHxw4CjAkUWkvkFrYXNEvZGK6bRUzcElb+cVHp86
/neBMYYcY8xWXr9OKxsiX4U9OgU4Iv0ok91WuXTkig3uxw8Wk4yVk1PS18sV1gloOu6w8xtwjhJn
IFLNsjXV3jYiqKwr01rZNJ5/3bRIAYy047aVUE/IHYe/e/M4SZq3u4nfc8on9wG0ekHl8i4dgJJH
8jY95qpEqNSlnVQbMT2GUASr2vlzQeRhZDA0gJvtNI7eUiluY40aGo5CaOLx2K4CFBZoLqHiCYa5
Pv4KFaHSDXNdF1ueTWUfnI8Iu0ObwTtC8UmiIVkIV1Ok0VzwIWVD7Ql+1Mr2vYBpoRhP/ZytL64+
bxl2zt86VND1ClGY7ap49VtHz5cXb4VO+4X33utLwj1NWbcoUniS+RKtT97FH1wEGrxM3E/NV35K
nC5aLW8JINKcP8sREPXx2oki8/tbn5PRdvoTOxkSUu5BXUlpginr//nQboCj0wJ6u60IJD0ABaV1
dscE09eILwQNglsiMc19k3MFINskslsZrLTcdE+D4B/AjcxNXXqJWXKDaqaMxYaPjD4ejVIL2kGS
FO8l8EDVqW7vhr3TmTKdIaKIKNJwkos+/+bdpU4njFuYIKHTmz9+294obF6HZtUEyDlZvNOXf70X
hirKhKu9NZB5KWgu9gq8dPssAVM0xa7AiTGJYeG5iuNP++zsumnbX3TXFKsZxfHot1o7y0ci2mcz
GH781cv7omITbxyC9e5uZlEFlTfVX0pp/0QrxQpAfRlKefHEGkHkqqw8vd38TKFsnU+ub+uYIhfn
rvnY9uEZQxm5OpdKds9LzpCZGBiheA6MJ+ot5tVBarb/6CuTMq/vhi36tMk5zS1eiGyOWVbqPiJw
JlBpa1cgjl+Lymqxaeoo871sQPy7GwbS3bvIsO1njyURbMwHHFuH3PpAgsZjVU4zxTDTWoJtN5jW
QWbT0XWNZrDuSfDD0D1r/AWpd4jCmoKHOtL6qp9Iw3xUVqjUbdJjxesPVNNyypWnTd5ACoSKST3r
g+bUAax4yVmPU9yPVHIu26UphOWG6ic9qMRxWkIqLooHprHbYoJbzewiyinfCy5UVDudZ5I7W1kx
RjDGFde3z38PUVtqSEsAlYqPXT8CngRXuBKVLZ+OeRWn8EwfcVl8ZWnCRv9FTeJ8wV/EwIaCja4I
eUQ5a1QXtq7po08ZDVgoPpL8H5CsX4jd8jk1prcWIZrLsCKL00ZN1JH10PcJEGz/fNqIRbW5WJkt
8Lwn++Bap5xNoEunmweOsEs0d/p8ncA6Hi8xUkpCGCQC+MMuMaHUxndycPJZTe2okBdNAY7xZ6+C
eiVR2fjEIYs0fRdwNtFJnWwfElmDl9IWBLbHsbFXQs8SRZ7LzGP1dVkDx2u2V13DSJb/z6zpXY/Z
2X6oLtIrB5k+t4jcQKAQogDQigxdepdZPaqr/wROroQyx9jSYa3v6NKz4l1jnrpyJPxLTu2a4lRo
Z02+YRt3ZEtfzAq7se9pif8tyAIR68eZpnYsi+cBY9yed/dSFtuCL144vQ1EICu4KRT1Zu4j/3aS
WmGx9kgo3yUVUf4EcDqsWrA3K+mNS32IbYHuvurxdCDchWwtZU4Hmp+NMANVR6zKkQKq2fQVJVGG
XwGOKu2i53a30RAzgz/uJA6v6xn1TKlK9MRZyqiS21AB97P6zzIiDR3IDChLYcR2/wFbk3iVdcyd
//Jm1ui2pqfJXTGXGHx+BB06OQ/EqoCrROgDLuflTYZZGPF4FncevO5b9XOrRvSEB/W+6RsoK3eI
69PAPlyii7CHNp+61jwfCF6b9AwYNvATj1T2g4SjyMUXDB8ggk5ZplZ9v/zTSPG1CufUX+BaUz/+
yjadw+ugY2TZIwlqE9UQkYmvUksKVm+AHCEh9gV5xd/xVWbDXV+NQSfPtudLkMSRBiCc3PmaDMiM
gSc6hwHEWeRaq6xyshsfYhKhQmhE8T3gIlZ1GOI4YZhtU/pn4Yoyat+ZzloQVjg2dlJ4IlJw6b8I
2SB7DlClsYjoJc/NPN8GvRLKFf0454K1E9IZL54EkIxnHVWXOZ5DDNLH/p5Eg4iIZNtOeEe1Ir9T
O7xiH1sxEtda0oLGieZZYb5uq9q/WzSBLAoqozQz1XBhPJLzNP6qFYyj/hlgYcnH6FclNmWLzcjj
VEj/utbvAvBCsAnT4XrXBo8GZIi7PVFIefCP41S71dj+wwkg2P95Tnk7zrhCjE+RuM6BCAwdh0dp
bxNrWQylwe/SpGV83aykRLH0NX2X5qwdwOyU+CjC2Whq2e85OwcyGcMDT8Mb8WWhrldnpj2TbCbV
0mZrwDf0z8L5MRlMNDU6ncH7yg9ZrIi0x2pNUt7qB3r8jinIMxDFSkZQaB5oITvYoNScozWnYMYN
NRth5Zb6fms1rsKn0tvKHrIjRmhF8IUdHxNqX2WWdC/Y8pqapk0wwF3/KqwNkqE+deIDCAaqIjns
ErY2NBpXkjWw2gb0uF8fnLXNcoTv3OioHcLlnBmelT0qZAb/iLh0R7KIvWu+bZ+EzX5wuIsStSCK
FrBRPnHMYhlkWdIqLphEA2WoKmFNQpzREKn9htLkNnW4WXmeFZutSjrg8wFzEQfseqbls1i0kEZI
4qfzlL7onCbfSyyyb0cHQVM3o48gBAewkhB0h6D7tUO5w2NqH91we/hBlrtdERZwdxEoaKui4nuZ
1kb+uS+7PPgR1SEPezT8BNFEQ+a2+F45RzcvMoWw0EXDVM+HQPJ4iCaPv/YP2i+aEnpP/SqyEkSk
Hs7U4I5AEsKGqRAlx6pnCv1pA23Ntk2tm0i8WBoSLVVUeA2EYSgPrLKTRvOIvHBcaK2MJB+LYmoW
HjRl7r48TdB8gshbTIKAXH4Yca42rsfLGGWI/c8SDJgchovbfxLHlzszV+zcTbCBcXQnJmnOF0J4
blErReAZ2WQWjSokg3NA4Ka0dAP6T6UO45HQBXJKvGByXMwhktp0aL0hyCBQoWEi2b4KkJxARq06
WaQYH0LH3PCVzrBPRZRqM5BSPv3KVsIlLlmiB7a5pCS+44QjkABjyF92Nnlfz7Nrr2Iuo0nZ0daa
3/T9Be7X9y2nv9K7bvbsTBNBR3dM88D46Spn3YpI390GwOfbR8FiFzuT49pSuO6ESEq9tnCUMDbC
J+0RVuTknmLJU4hhCaOa+fgmCBZnl1izO61mVCLYPz5/ZexBhBLykMOVJQmDC0/B3iRu16HaK6dL
3R2oKtYrbvxMDNqFt0TuaJAooGlPg/tm0nXRhNI+LrqAY/iKqieN3XMZ1ujdUQnK/6vTRooa6eE2
bw3vZRX7LDS/+ef9iYaSi26M3Vfhkp9a5PSdC0j1Rw7AQ/0TmoTvNlYiGv38tDTkqkBmxspAshKV
TSUZTaQgefWsIsKQxxbEqtpE5NYav/u0vSfP8iV0loDSeMwDrOu+4m5YaElX7cDDd81ZqZrYkxZX
ShXtJsLElix1vJwdxfyXlMwNrAWslwec4DThUd05tjF08CU9QMPiQBzT97hGl1RTk3zRONKk+Sxb
+UFHMzKWI7ZKbRQ138igrUhYnqRYyVTOFTtLR+kCCsJx0e6aoRUSnw2LUaj10mTm0hKgoOeMJlFM
G81rJDJnRIW/8WG/U2hjbZzZW9xPWXRNXGaMO2XhdLKBP3u1RloxL2H8ry6jjhiQIbx4ajCaCWJm
XFVk/Rbqios7ZlItuhNTiUfDutWykeU54luAmV1/9EIn8UlrWo93CH6deUHho/xBnTLdKpPuy7Eq
EWbuvBQvGZCLQuT6dO+KYpkJythjXPJtQLwTLWvMjTu/cFCuEdtWwDJn/C9FOcTVFQN/jGg+ADLN
l3vINgGufZxwVoF6vaVJo9hFnIX+zygku5e3UmIC7CdBs/gfFOHKqpy7Z1HrHA5Si/YI50GDG6gg
ky3bQBOIrIaEGR3qzs9xnJAZzEjKTAb9ekWoRYcgeIvm49c0+6kjs3Zmy93ePM2ks4KvsG40gatV
7cLIUoke7yfkpJbztiT+QBFO/qyXRwtkGgVh0u6+MtJTlzoN5ufO329MSS9FAVgDC5/+Byf0uEKy
LIRId1wHf8SqUHhyElXGDI6h4gE0Cjsnuni2HnifUrA3PAzaoDFEK+mZUESQeXYGiijujcAqeAa5
5QGTa9DW36gN5G5BK7+QwqVJ7sI5NQQzdX33NdpzQXHzh0eKSsNX+4EKQODtSrdo4SRjAe6+T2SE
NA1XYHfj1WdF1tqxF9Og97c86AxolWm3tvkbVXpoa1CNwjFitwzmteI86801DB84j/N3wv/wBPMv
GNDzxd7en4Byk834mvdKidT3FYfdrL/gHVrgTRwLjcv/Sc/o8a3yCAVEQ6wCtzZzpgJMxrjgrcFs
QUTPESm2QxOqvP7+t5S/I6k1P4gEptdIIXMBysJ01smET8YTm7JOdrC9xASX+hg4U5nFbxtmHXSB
ZOjtVD7kBYqYU+793lmTSiPmazcX5bOIK85tOHEPlCwOrR9YlLyQd11qOi3fAiN/ptLobLhM53tw
y4q2KEDuuuNaeTVB5Ro0VRAverTmV3PXghYMkiNMfqdEVr64hOIMF3qQrr2HzNP8OPz0E6q+XefI
oSeM9zA/oid2jdndKmyump857vvM8mW4mqIh7jIu8u2r62Kp9h8b5A4aVT8RoAUgGc4i7mDEHGLO
D5avpBwTzgfO86YayhxpnHwG8yNyOjXF2ecmrd8cOfTBM3DMspl3MhOT8AQm4V0XbDen6NB3SDNx
KpTTnDNKplYnItjrTRAKVszQ326zgmtmmoyGg9//qycNy2CuMU3Nr3lUBPOtGFBE0RldCGIPqooD
aoCt32IarG4HSbWlTA78Dh4OHU2UDr3QXBxLt6fyj4pQtsXCQvCfyvEY8BpOjEsUAysSm9s0xaqN
I6sJ1A908K+PYLbEKSxx/gvuY+T02Elmj4KPQn31FHOWDLHrJqh56CS7U6g1nFOn4UcZ7HWq7khX
nE08vv2wanij0dMMwY3yhLZXv/i2HKkAnwyLtHpQ6bh8G9lost5Wh48TlcwAI51MgyIN0PPo+bfQ
lSOQI2jtqk3GJtGrmHIVoZd8XVozZcRNG0TANuQNLTwFAhN/6MBY3Sx53BBhwzt0Qu4UbMHnjVSI
nAstjXAwpZgK6V6LIELVwg1rX8stxHr1XlyE4qsEbfpeqNWwk9fZgpl8joI6wau3XI6ji9u8GVfa
vi4HwVIwYNU/YwOLPyPBLCZBFB9MSq4ACY74nMoWgpEGEexzBxfOVvlkeE1UiT0tvw/IiRmLgYmv
zpZnKYXwSu5UNGk9Ld+/ZbTtuHccIIKkrWp7AoTDO03Vv6/jqHh94a05EtL9uFl+/H6/lP7UUdpz
dIALJUOTCDV65V6w95SrTJVpy574hQEpCx5b+vypBxfOkMPAtklqx96rizyBZMpAj6Jd55YXX7WM
51bD9drbxTCxs9qAmJQA5PgVw4lY324nEq7zsGPtUMkKNbdL8KannuG5Ppc/Csx9BzTdWG89t53P
V/Uc0wkVjTpoToLrs0ZvDOraDuh2+Xkhhb79xS0tX3czvwY6mJNSQzlYo02vbmwS5dAyxYz5EkJi
t0W82JK5mAQ6iDN6Jhmx7C7ZUWGkYk/UpsZ9jKR5bH9eVa3g6OwpbUxtm4aSu7ZVI10NOmzwlypI
IRKq/PF4eyTejfLoIrf5zD+msxefSiOc7egheLRGT2xW5jvL06FRyrBmf4WWDHl3JFTGzeW2Y+W2
M8CmrXDBGYj/4ejl56dh/WYMyy8GhorRWGcxO9O5RKK1Pfnur45ObtV2pwrgUSGEtETV0U/SQa5n
LrrQvc9kcANmXpHaSsHYnEsZFCenLdGWEdwXFR07U3j1ino7KyZfMrErfOs5qkTIkMMukAxqqz3Q
ADTYtv6ZPazrN+SUNrhqgQ054bGzLNP2tZ0HhwSd5QFxhsvKa1f9YMNfkqy7wLDdZCyF8BH9+r2v
6CYvNg+yVR07y4YoJt4tbzeJh8WVR7V8KSb4mQZSQ323Yok2C+EYtPwSTYFFid5D2DCawc3ZZz7r
HNfuzeYNVPXVgBYKSreRfh+D3BRRjSiludKy1Lben8SgK60B35jSUcA0GJAtYvK0CmIRV+PP57aV
qI2+ArRgXJpn6novl0UWSbllA5DuJcF40wa3gmGA4borirLM8t66sPB/dvKc/78SisdyS7wfsd3M
lonwJtU1dXUZe2zvO0nqe2R3E6/h5CU3jzKnrf3AA16Vj8iw3QLi08IRtB6K0Woh65hCLDd1OfJT
aqpSG0U9Kv1kRBOCtM0oLhQx7BEza2n2iovnd5ux7GIMFEbxD5eXHWPJo2+07H5yxqtsY06mXPrg
hb4Yg5q+KkBzU2W88wMZXwYP3W+0W0rjQPCIS0U4+d4Tjuy/EwEhj0C6faYgM3tjm6NuA/U396LN
M0QutM+7KHhrnwLdxIfeROuPMSP7YDsSb8wfyWkaEemoSiTIA2P/sHeWmZ64hmwaYAg6P5tTcC5S
vECJ/F8wpkMh66QvwJncFXBI2ZZcgH7fUEbLz6pj/3+UbkC5U5H2PEYJE4ZdEdwezW7DEYivn/I5
H01h+TCOFKtw73ExptBrHZU2aAg9Eh6pCKHaKbWJ9V6sdxhULWxGXfQmFd25vL8vJWzorCJk7KZ1
yb2Ucbbd5bDalRJOPAgL8bpL+WdZpQER5zu7fBBkX+77r+VlQqGCemXkbaJmju+Bv/knk3BcnEe9
u3Nk/YAyQ7OmJJv7Ze/xWCFrxd7O5M1CXykxJk3oKaDjBv6So306n+dI/71B+3N3p+1VS6Sm00fl
QlWISTl8A/nvydaayOyAVNk80JegbWexrzkywRexiPRYZuxhCT2E56ugxFjLeDxnlpyUokxkTDLN
EBXI3TODpHq31TIWj4Bb9uqY/xyGl2Q8H99w8K4W9vDM3xy4ndsKFmH3/aRlaM0/2btdrAQQhDXw
Wq+PeejQC5o6H36U+5o+VADGU2/+kpoaq+Z3HSsA7WrpjEG+4RiEb3ki3STlOVvxhJehmkQOzG91
2DbG7dBO/SO6IjmDzekziZM9mLWH+ZYPF32tPYnAaoGaZTunGAEC3igwdLkClJ/6uHk0bzJSPhIp
QsIL98RU+P3IuFOnShoSRkb2rrSa8a1dmtZjZKHMo7nyAK2hHmy+v9wffrohvRnPSef2evz4MiNn
p3T0lgMPeceyn/ny+elLYEbPs3W6ZM2agJCo/Y9ib1NKX5U+X6B3JBQ81rO9mt8NmqmpMoVB8+hR
w8ZxxjzHMwLeoFh0F8blxW2duIlfRhhZBLnqgedG+Ku53BRB3XxNtqy0TfnmeX4xQgL90tKAatd+
Ap48QA5dpoEcx6OztnQUWw6i8hrz6UpOcPRP0cWj7/Zk9bQUGVHozHWzBPUZSY0fux8cAG6nGfMe
pZNF1taakeb8Z8SqEnP7sB1DoK40bJI1ZMs/VXhYTEhrj9talNbmsq5Y+4VCZs2NBbDuZQJGMfJt
7qwsoO/aCBAXG3On6fqDU/XLa4h30OHlopUaO/S7Kz5MavHsq+l6KhA30pmABD094outJILEst0K
jNUS9mj41KSXWoZexvFw78N+Ueo3f0DrrWVxNA4QMtt5T1YmXKI9DQ3ZcFLxVtMHU8AL+R1vfoXy
yeQYLCsmW8w55YCUjRyfI6Z7T7R+MtI06iIRMBpk1RVTyoZ7xw7VXDJzlyj5qJ2j2MbfFRyuTjrZ
we2b/AyjqkMQWexSCqm6Ps/XttQ36iPlpAfGKQNEutok8DG/adt9nziQlY5MMpL9yDu8pPCKSUwy
YU8VwkuupyA35Dh+npWGOs+fl2Um27xUvvuDKcitIkCLK8lpfFZDp81/JPsnwoAFmIqGjbluj1TJ
xXDbgjOiO2AYPg8Kkme5DUWF3PFdOcdPoh+Wd0tpXfpKy64dYKdOnxa/B2haSo7tZ/84eJy6YpEv
BIiPfEFEAO02O4Tqk8pBdF2lTKM4YaJfrViZBEnm3cUU6c8J804lLAjsWEoAOQ78SlNBu0ov8uw4
2gL+J8UuyzHFKeofAL2szLsgl+s3bBx0IfkQ8bPzgfWVYEOGJg54z3KqH+Rz97dyLqfqYZHvhbmv
qo7Q62Q7pFTE2xrZusV7qaKWZR+Eg46lVk5LbMJuCTpMKSfPRzpUV0YxEf9EJn7sTCwtO4HE+2yJ
yZGsF9+ViHRgLbegjfEGfF3WmNqMUDoq3AuD2A6YaB67vJCKQgwkW4elWKK7V1dTs+8aacUTbyHq
5HE9v6QxFJfFYX+u8TvzVUI5hjYuplVgRCANwWjTEo0AXSS/r4B1YkkJoNuSP5ObzBsuMRLuPlOC
eqEQCTYhPe5TJ89a41AMp3huwj3G1e6HdlKdQpY6dx8aSL+C0mMKn/dY6yh5gHvoJRLooAM6Ovz3
X4ASc3yXf5oXgAcRPzZnimcO7PvDwciWtC+Ypbi7ZqI7MFxOo9JmVxTqXdFFBpW6QePejhOfADKg
lZmDgMgWtUYT8EUUeMDx7E26wOGPb6/CKahJtyxdso4EOBeF1le/m94Ut42VwaPVauG/E20AFTOu
H5uScxWl5Ae2ficSuIdVnMOTzG86k1sDA+DpIRCtIB23zBZUusM7MSzykQON7zDvirSb1p+pqNGp
ZxbMMlMVRa6cIM4oX+fk7NPIA9GghFsGYU/u4hFqotjG/F7xdM+DAfhLzix6Y47tKRoHjeByY+Dp
YKOcxetDwZ1PhIV861pEvL+ytjHXx/l0ZeUnK+GIwtNzH6Yyjxam4E5l9trlzNqk5GxpRG6rQEx3
LG4fxbuszHPCvVxJPgj/UnzcBJQkNqyCNbAiOOUW7Ui2jug/iWggoIOKhYeQfn9g48z5SstKKdoy
qiqat1HK+PNmA/kMykvWYK9B3OIv0ZayBuyaGxlgqJ+EmxFKvba5FTXY21AhlN9ma/pbDoYH6mUs
X7Dfpw6EOavczKo9iv1VuCI7H6RNnztBRnUR+Y3zWvUQwRhOUjengo09bo+F6LxkKLADh/sfZQSz
0UacLigb2HYyANj2WFqEz6d9vNBaXSe976C1LlEbRUnjl5mM0Mfl+GQW7m5GO2qszRINPF8L0aDZ
bB2xVFPT/proB0vQW2HVKXK7GTnGOu/lN+p236EuLhwe4/Bj3WfnxWJ1FYhbet7R3t4oQ8hXQ5Z2
Pa/zBw6d/27zEXcTnh1rtdANdHkGHBpca2NQJ8Y1QvM6XEoBvXuQyBfHntKIxQzh8qCSj2W1Vq4w
8d3uAe+qlicaIO+V9VwL2e2CeJaz1qYNTnHflQ0lsbmgK2zKnGjGVPvqSlWcTjnn9xry+BPmuYft
FF6rsFrnc0voykV05eP4S/LQVAR+oFUJaXsRtRil8bSS7GO2habJhGIr3CKHLPlltEk+hX00vg/Y
kIvrpHOkqzzOslWq86QD/MAPGyEFCTfCJGH/xKW+pE1sqTijZsgO7iyf7/3Iq8O4w4Yh9dh8nl9b
LLkdsnMLu6vkFIn9Ny7BdRgfrZaahiIhlVOGppM4WJbJLRL1TrbZJoOxKiNrOBLlf+G52zFkf8ZC
4divtC6A7jTSSoMWiE/HpPSU8kTxzEeKJXEwNdtA1SB0JYr/AuSAH2hB037j+FriqYzbUcDkD+lu
foh1R/PciD9IcAl2/u/GoMm07RUd28DBcchImg20wjfNQu3EmPo1W/66rl9b1qPp38alQIaegpB9
AF2VrwkjoyCZKYymEjckNEW/XGbJzPGlf2cM8ZCu2mTEVr5bjm0el/3iMXvJJMjZEhkO2qCC8Iqc
t+9QmsIa/1Lr80ZBEntcoJA4D+bueMgx+7mM8EnwSUX/wyDJNfNmXhmSnq3aN1ODuL/JXlYOUP/j
o1vXR5QFzK/WLAgVm1ow+nkgFVBv1uGDUKFBPosjSLIF2AMyyKtAV5qwbA/3X5q7bNdKvICa5KKb
6eCMWsiSJhf7sLXqqGuB/fMljm96TSnK4ntz6yc+5WHxMVXqQLI0OnhnZilioh/8sFvZwCIV0/1T
yTLzooai0erdko/Q+7H9Ky7QMcMx/ZUDIHviXFQoJu7EZMfKEDorpaqSa3F1ghViYjWYgcA0ZVq8
+mj1pzpSN6rfo+xNeb9qHpLi22KuEOIyi0pARn/KLeX4JAlZFdXETFAUMrMEWppf8RV5tWD8WlGL
TYvVXh3E3kwsf2+q9gYCj/s6lLAfYjzZrXUoeQ7DZnKpNVjjwZX8Eml/idprDcG6ARDeICl6Kk3Y
SMik0MlRWDNhAH2vTbEm6Ut6zXTiiFMBz7xMaitS2Tq7ApcuQnsQJs2mwPmZNgKh7sv90Cg816ru
E6uOhUeGFwoIUagopuRQfTATmD5fNTGnt5ASTB8J8PQgrxDGSwpfWCIOxPIFcXX0BudlZ549o9o2
PTsbk2Wq2WsbbyiOdKOiHv+bKIhynwsW9tKXDwyeINpGSErzz/0MYIvng/GPQWoDu3znxa1LvY0P
OgvOB0hzIJgpj9DEPZ9w4bEVM9lWJjVneieYNcO/hq0CYK+ZfSM6I/ltE4IShicDXS6TpOXP1hB2
aMaY2Qgp5b0DH/Emf+FUtbzoagYQQ4yjO0EEKNRaOXG+Elm23dKuDKjEH8dxJzJ3ZIpkhMdLH3BL
kY/2zwW6yrINiYs5OofVBORp9QWK7X95Q9n7Qt0j9cQbnWWzf4neRHz256vFx/bu4q6EYhhsxaHt
RgtjdMJkd9EnjGJ+cHJPD5uNY0XcXWG/XdJY8MDKRzzuyhpoc2/ZQOePfEH16EgOqf9H9moa52xf
MQduNdO5/eKJ2lHowDJ3HwPApj9ZfM7ahf+fu2PZXR3Zke2WxNMoTcMMo3eeDD7u+ba6AC1FmiIH
mHw0tTdWNPR79s/KYFHneGg+LyMwDkGYETagG8UY8o/1iwqUJYRwByQA7SWoJkF+DfjfZlVJFThy
tCD02vaXv/4nEOTpUYgTEEYABkG0uRO2U4LCrC66wSy737CAHBkDs+fPK7k3t6tnnK47hmYd/mQZ
RMoO+YvO1cJuy6tokkGfyNutpLspEsjf21PfzQ1LnjIHwJGYorsTMb97fxjDcj/C3XrA94IgXGKK
3cCrYQRKqV4sojxNmwHyr6OKAhdbs6iX2xMgn7uWS7sBnC+qGrrL8A0a/ul+LthUdUQtlKF0QSfd
dwPCybP79/+/jyHW0Tv6UpkfXhQFC/1UOvqADhBHld+AZkkaiGUFHgpbWof0PVIHePdhZ3F69+az
1bmgyOZXSLQ+RQ8xgGECED4RXIqk/L06v6p2O0V90CioOBzMhqjpWJoyf80ra+XTPC3k5Nf0WNAE
YudLKgfFnqtffICB0WBgvj1sW/twR2QdevCTeeLj8PtjNUA77eIGVhkpAtOAkaf50vj3R5jveAj+
1A042k61nUYFzhVvzZt0EBC3ZnzN+8R0qL/pFbGcTKOQxrM2Y+zKAfqzeoXb+GzA0YfyRMX9VIbq
Q3eoaHra5NxWvHn+4EtZuRHm77bGNgOXaq1UlPJ5bTAeYPJp6zjKtI9uZj697tDjmi2IcgLtcM8H
ZZFoPgsPdFfTATwaBObV531khmhPselyr5kD8NHk6rhtX8fNZdATtiiiQuNGh3LrnDqgI49YUOX7
fpIw5W9xKCtmY0M1ZnfzHq6ogOqR6WE7/70JqtmLp2guVtPtddPgbzhsxMKKxLJx4U4l3uYjuEhn
pq5CDWWxUHDMhPN8swHGWlz4fis/pj+YMWtzKpYs9vkgzQg3Ptb7YfUc35HnxAMfVKEbFiritd7/
yw1AkrXlUIyzv545JBJIXZQPXSOtsdr4Hqk28iVsAR0umkJ955vfmCQcj1FUtcG6igu2OK5khmaZ
V7QomXGGPhROYINUMMYNzxZhOJjoS6APJgjBikykbwCrKuNy4UUStkcAJbi1En48/WlZQulF7tHY
vtkj/zwuS9TePLSVMN/LYx882FdE1ACvnaXYZOKqfvJvUbzRE2FgNLwzAYkzQZG34+COVpq5ZV8h
hL7o9UP5vtPDic+3fXl8/jdBqEkdWEA2ppma+SrXBaPuf2AHfEtghuNQe3WBT7zXFRTaREfxCoWY
LmCZUULlueQ9MkjlIwoaed28f9qc1PTph6fzeqsH8f3HdaIg1e7MdkUwpSMgfQx+BJ5SM9TFwkMA
YIygjeo3FfdtLV0oAxRaJMGIsxj9brY1vT2MJNvO/oI0GiJPFGOKV54tGRdr2G1H4oywcuK/JpjR
VxWYc8El3dWBIAl5va3+pPdqsXvtA48XhRlcMdhK3BOuvjmmdjNB3l+s0BLFl2tbHfjJL7ewJAP8
NXqL2FX2rc6XFgLLcdl6e8hbb4rf3vVCPEkkGpvKnTDI7qq4tX/wantiQpX1PoNrRGCNET801Un8
/bFCF+spROH802RB3OFCLSEaoOiq2yLIl1G+AtYfytvSTL5VF2r46MmB7LCGntZFA+bMWPmCQngD
wFJMmilsXrspEkyluUf0GJjYpJ2WfZtAmaSAhgxriC0CqmT/daN4mcDIQ/u2HrfI2JBX62IIf4Ad
9EPsA0M+fRTgOqFvWslC4K2TnBZaiBxfgz1MufboKpOdrX9l286BROKv11I4/hQsDiyX1y5W5KM0
K4Jh34BACNIggunYRkp/8cdC85dLcSVbWWRIFppGLdMqBdX7g/WraeyWFgSY9MDV0kfygssacBa+
dxIz72eLGvdJw3qqKh9SUGT1wye+eyFybEVVDq4FZXEzP5q3rEKjzJth+HWPb46q+GeVYF1i3vy4
YWdYazCePAQ6XYwAmWfKylkhlkSxE805yyrnneC0HXHfu/D2TUHPHbuVtXxTF+zpsgAFzPE5FEsf
NGP1AZq0R2KzPQU7kTmsNvEeLdAjnGrdEX0DEAkKB+JgZdj+z3+AcIUs6mcYKTVWnMYz6U0T47ec
AdJNjAqNapEJNuILMyRIqzz1Rg+EhaTwMsxK/khiJBtGAZ7ktff+X8V7YJJQbBkMNbBYe1y2pqWq
udQ9vS4EEMRBNexvvBnjyTbiu5I+H8aFVgpLK+QSe+Np18C6Ezvhu5pO1i54TnvKgV44vFX3KcYh
ML0dY/2nEtnxgmEdNS2td1Jhh+eQkjwf/iWpgeaBjw7ovQUmUZVLZvk9wETvc7fBkwmcZlOY9Skt
EDQ0MJ+3RrBuFSxsIaYOIR1GqsjS5Y5hn/8A0vye1/0jfUPf0Cb66GxIgQlVFS6feHbvyRMeonPM
M0uChjfsf5XRaPc9VWKPUZovYJQhNfD4KBMegMI6i9GrXHa06wjPtG/rH5UEuKvXUsCrqxKplMVp
2b0a3U9b5YKxJEVMXeF0EKqSC+D8fX4sx3Yq+wMg0M+Gfn/TXb4sZc8YPc1c1NsQ+O8ROoI+Qjaa
3eCvmB15DKaQVn/WHd1lw2sO2s8/gy5OUxvxYZXvtRLDPnW1OdRQmqDOPL0RqoIfpCXOpuFaR0U3
3+pOHnLYn1/oRkyWeXgF2cKIGGMrSmnIz8laIUaofJ1uc9aW3SfJ6/LtJHxZUjA4sAcl4XNtUV2P
sKevghJ6Ih5Tc3s/fjQZrJQziGWhy6hnS2Z9z5EvNk0+hD5HdmuzFVX3ip44SpD/fKaM9OV3WBT4
ib3NGFBOcdqCzS7VsPmI0PsbQWC7PYFhHQ+27PWHnA/X4+zaYMFA1sArsSJZZXX5R6Yyhk4bihFu
poMLT06DUZvATb3onEw628C1oPcOsuxMHL41JkVO08It+Sw2+YAVNChkfbfrF6P8djolzy8j7w6r
+dxfA3G0u9TLwEz15V+pQqLM2mERDrN4x7JvMPO9+KP5Be2riuagP9mfsAcW10+KQqvcNBLXvJDL
V4Hr1pZCnUmjGTobw2qKuBW8lYevkOnGua/oPXhhCFm5eurQfsf076eEgydUU6H6RKycLmPwJCtL
oMsL/YzcwpFYh2xiVsWzXPGx9m8yokwd1Ol+j/y+I2eJFNbdXONL4GjTxEW2XyvXAG/BePUM5bIK
HxV1jno9FKqgg9aoh+jpOa97ZvaNtWHzSmXZ04jfLJXxjBAzk8MLPqNhzbIB/kUx6HzdZR7Txv5F
KuWDWAgQ+1lpBh64/TgPIL86a76ucKUr+LoMJeQtZK/ce1PA4Pji9wOdZVD8XMAg+tybbdtcjNYx
1hg6vuAJgaSTXCNSFfkXDqx1Pgf+LCRfujpdbPry6K3o1FZuNUR8imCSWZRCBIXcWsXjF2mHwzz7
OqfjxHwEN2hRh9qRJVWwIADM9vEvDN9ULixmIxZJCtok8LS8MpM1HxZt5nhOZ94DdUmbWw8+61RK
6HtT1B2iW9Hdz5hgQT0A29Op/xyY4t6iGNhBfPpvd9v5Quid8rcKYqFv8onen5dPUwvY3B9qX50J
5OywO2BjytKfCDCNi8J3YLT2WErwB3dRvxh8BbLLVOWWJNykfJJ2nw2hdS2MkZ1Q4B5lNLBVQI/j
sWnFm0sbPlM9mPMZ3vDra3wHPvn3H2WmaTaNzbbCF7p4SjV1a4lcfbSO7mctkbTk5l2mibngYnaw
kn9dTzV1eWrix9ZbOPRY5CjAkR4Gzii5GVINsA9twN/ecUSjymE3deY0CS9dZqBslK2hyNwThosu
i/UlqJ02tIs4ftCeW7k+oTGIkCspnr65EbS5hZXx/uPX8FlBOKbR3eurE0v9vzt1ntCE+VNQYeKM
gdrSRheLcQBJswoY2OPKguh57IL3qbCjv23TQ1YIugjwuuBgKt771VKES1ggA6K32C6pGwqxSWZf
pkoGpb/hfIhi8d6cKldmbl7ecaejYnD3vDJsY+H4yKZ2A9hWCBjD+XQxA7UXUxZmEy1BNMDipmZj
xTStv7+miBFI7Mv4ymOCkmXLR7pDsRURBTHKDpx9Qd1z82OCQ9WwuOmYzPDWJw/b5qWzjwvTc2ph
Hhb5RNhfb4pN9yHr9jUhUbr2+wwAoT8wD+ZbouLXSnsTTXwO7gGFtiUzNMO6+3qnEJD8/i7erYnN
Ife2TZTTEwohup1RzZq2pLXVtYPHHycfUyD5YJIS88EonnN87BpWzyK20ey1KJumC9W+tTz8CMpR
mLTq1theXDKbNZAKXAIFxu8TMWXaLNbGu7y2yF5E0CvywyqcoUONFlTmBO46EzJAe9QhxYjfrgtu
cYzC/9M4KXNftqzZa0ICRy38FmoxeoNqelIDQWP9LN4UA3YEk4KYzduBRIZx9oFgolhmnBCeRmGx
KLambjC5K4p5HOGYQ00cVF0BZNh+XQafqhi0bXjr7QN9sTUX9yUfGq/qOi0Jn+FYuEI27Q72+zsi
Hl1TfYVKzxFerkhtdbtSqH2rnY9mqaffkl/pgftXxVAO41JvlDeMzewsOuhRDU3t8IF4f5BBirU6
Ovqr9rgPSgVqe6Yi5umtpCebiYkxWkVZgSiiAEqbRZ3LG/8CCX8fqZlRQZcKGyQkQLPVRtijaJkp
Yiiha8bFqaSWHZkSiCYXScLKY9M7Yhe21Lcsw7rF02LvP0hprYu1948XYUMBNLFkc5+28LRoJslR
hThtMgCroqbcxUHbiKr0S9DiXoINR5j4XPwLNI3De1dplf83tYmNxQty4SeJo/B3fIz8jMlGp9Vv
igFjb2h1TurUbsqd/fDC+8Dz0o3cBDvl23BJlY1uBB4asBBddvSOHv7UfdLcG11l/IomxuCHz1qC
h2d798wHPDLPHnGXy7/wWgXPM6FCPwjoQXsNpiDtmizxETM7AnQomQ2RhK0U2jBJpC1oeEM00gmh
D4Ws15satMwRyqHO4ZiFNxHeOVhwOpXdDCWS3QoLUFsIMGGExTvXhGOhuYeNV5GVi9R3Oh5n7flU
ykbSJreMZMp5KPHPNs2KiqMAaYgw8Lz9xNZkB5bd3BAwNUYlzvMf7SNNKvHxMXifGL+2sHRjIrPL
LGrxQ0GSGbAvhEu8BxSSYpHg4lZChkzGPeVirWgE8n88S6wkmTvXvxsUGGalir5KXg6ExAjQy9FU
kTrTQls2EUV2I3+Tv4BEm3SGcJljTP6n6NEsS3530aFKQySv1Kq5RlVov8UxteNUn90BwTnlNd4D
b0M/4i3PknVwi7lgZMhYweZHhjgDdd4kqMFVbdyCKfr7n7V3SBP34UueD521z5E0iZnTJUXpYms1
ALZYLe5HDSbHgUVLNFCa+qZ0jgsHO8iZHyUuE5xNezxjeNsW6nuCxniT9tbto7sLWnQYcT5Gst5z
SgAF7LyyUPu+r38URe8B99HQAb1rQpvOr/bmFdJge9M6Ol9tdOKdAUdU/5yvPtxQolX80CXyomsR
SJ+Yndsu75CADbmyfoL3gw9GAbuXLdr2Vq958sehzQO5yk+fkEVT+nZUNpDnXW7urqe5dg0HihGT
TQVxiPWy37xGpdVOOE7KsRdn5XAvjDMxhOtM+06u1BVWTGDXlp61kTDwxjFomSd7sAyWSchrOqWY
/4gIzG9Ez4pqfsXw6AqLnk+paHNgGesi3jUKcbigqpZzzCYAxp7NlbXWSf3nhqT3aUrXa/gY7i3u
EAidBYsrGhCg9sBZpDDj13BhT6Bj/lFT0CVUfefiJzt4dORF5Yg1vJmeD1o/Rn1efcGChORo4R8w
aWMozLgPdjuYy41Q+5sgFk3XLXI8l5cN98lLdOGghTD/VSBEMipah5HDIqsms5tzJ67XeE4s+vi1
2Hkadx6oOY26gnbayFuavpyR0doAszFhA4ICGJR7S1FHqtVhahV8ODNuRlNxh8E5cnkSxSsKPiDt
6MB+cy7G3TujgZSuoDHOhTmcBB9GJ8PRp0OgrqxAbJZ2auVcQeawu94jXq7IsaOS4GQLuSK/Mg85
UX3JjuPO9KxmhT9qmGsvwPf/nuiTviUgBzW2iJ+msDliT9H0JF1rE9sWd6h01OPxBaRmVQ9pnhXo
OXaT8F3/wfRF2s8gb1m1HuS07Edhk/uNyYgp0SAnGyS5wPYX55Y+bLn+B+mlwbhmvFLpdlTxc2rV
whLF8wl/XppY+i2UvkiG2Hz7i3Ifl6StBPzCEEG7E74ZJ0nLRNFDpnUMXTIpTPWaOKnvAvWpTn/g
5VAfevXfrunfVViiRsWixPqaCT1stW0h9c/dCE93efQaK5UnTTbg7Rs6Ho/5yThQtrBrrKwqPqbm
FxivlRMqmsdiEVUPs0lVbPyPj+ItI0UrU4eoZkWUcxK7V6iz26+NykyO3iL/NbXbLkIDZWtwwv/m
/kMZbentnJoH4g31HxarvE4xCjG/inAzc8b45EQGDoUfbXAf0P91+K7UToJ5DNq6CxSUFj+9hXQq
BfpDmJ5kHd6Q+AlAkCxROHwKkibYptZgt//UyX7eocjJF2xoP2dPyYLsBaUBube0xxIDyeDq7s60
qMxqya+x3umblbB+4bWoRMgdNpVWC/uTs0MePbEmFZWARzico9VIVqcgWjZeKZNvgkLS4rURlaUq
s5OFNvkk5yN7qych6CtvZncBZP7/mJnQVA9Wm8VbYIiN+jPxGtgPUNlmULHo9cAgu5sxexeI5GPP
JckA9Nc0qLwj4ozrd/+RxRrwez+msiBWed7x2xCT8DuoUM/ixqhLZJtYp6h+hnRMt0zR6t/hSNbA
n1jaBgCMrLMl0WmsgYsBuYyI16czt9yS/VjxHX+t1LDgGEIkAnIJtSNuIUKr9n3My9sd+q9YRCH0
8KiUK0bxnCXWr8TDHA77/1X0NtKbHIl4bJ4gLFFZPT48dwa7D6fVa3SscMf+MDHZ70NS1aIXw+nR
CevpF/CADTecp1bQsEvT3arAcIg7DEA4k5VjS199CsL1p7/FAGhpMrveRlQPdj9bMPkiCqBKhJtr
CCQovXxLJ0dk3N/i9lqRhJV58lKzhjgUpkxuX2OYXtjWtBOXxanUhOOHzLQ8CZYNBGLzbBxeoLOC
y7GzrOCDrExOciebF0HfYn+JPlMcftJs7HmDSohwhoJXSLe7bVkiWNLOGWLkzMAjxfhFLe/tNWE9
c2eZC19WvQsZGq19GRgCk4PDT14SxoAk8HZsxzn8ILHt5hTc6oEdVVMM/NMpJfWb1G6Sx1l7usy5
vfqmwOrBsk8VPB1CFNPW4SZ74rJWZHILUUL67F5HF2DJDGj4TEGtU+TBgZzqgIQCv8zyf2gOPISn
ni0jbScGgymJLTAofRn4U09Dyzc9pClEVg3Oz9ES1lEXLhlzBe8ptbrdZJs7H0YF+sW1khpDWrkw
EykqlfrzqO/LV/dl2+I0EOXTU6erQZUw1XpSGiv86vDl01K5PFipCKvUeBDycB5W+Z/eGQBu6Psl
FUAST9egh7+kl7vrhtSzbMpy7XAo5ZQugCtdajyGxHZ/02CwCpmM/+iqnkbvSpVtdOp2U4okK/lY
haVjcOHlau+HU0p9x8DzGp6KMQekNtF7B2Q0Od1s1qSypiB6Y0EVcH+xL/8f6t1PLe1cDURJN2ti
Iz8fsr50aDj4iTbiTJXgNWrhfcPPG3fjPqIoaSs4ajGOWo3GDc/u4C8wGCG6n3zCiioMGhoQJTOD
tjZUF4DXJzS/71xO0XbRLjSDKPs3R5daaKPVtfnyBBm3N9QJwQ1CBiJ8dCV2QSk6PAd+6FUTmssE
tDiWiz2XrLiSlPpdUuIc1/qUriTRF/MYtqIjOa8BR8w5H8Tz573vPZC7SUCMTcZ8x1tC7dHGAiCe
5BGbXuIvPX4SQL+Jpi+f6YqquqpIaTdod98qyXsq7H1wVQLwI1o6lsYZxNRFYj06Lm7A56SqFsXg
nFNObnY/IOFT5L1QhOiDyElwV4CZOk2IccitUijw6AdrxR9jS686j2D6sJdZ3j002icngGA11Hw5
RIiGdp3Gno/ZYW0PIXbDvFr9y+JlzcI6OcqJrp7/CLrjpn8BQxCFk8wQpboIgtMxvMDHeEmz/zjC
t8cHle6Coqe51BoMYwfhLUiwxvaSWl9mg1nOptJCmgxG5ZdFfUHQV9epXyqPF3CJKke5swF507tQ
cAjMjygD1hSeQtf74zv0g4oEYS7dE8EyR1yvs4GMhcNSEtqFU+Yyev2ChTBbCQTZNFLPg9zcg5vf
l356AvroDrZNsXDfBjikQVm6KIyYTmoI5svI4j9hiJ6/reR0IGVHikWZ/78yYEKZpfCewlSV2+FQ
9uL/ZUIDU4LJg0HqN/QFO4mID6/lc8a0OAp12f8vo2i+dDlfnliAPtGQju6ak+MX/woOv+vdXRW9
OhHXzxB9TaxayIHw5ulCEf62gzAWJF1uzqElarzZEsVy/98awLxaFxNU9GJzOeX0s/dcvRdt0YgD
smlHdCSUvyHY5Q12Cabq0HWQLkSOsVD1h7vWOAq0RZwxUYTJ98sfex+DtSNhld4r2EC/3qSigPmO
1YVT1tSVXmRFsqPm7c+7W2GnFa/jfCWFrPST2dl/0UBflgIIhF6vGlIq2K/ragLw6Uiw2FiFVD5K
fU//RxP8u1edRix/4EorqC5j2ZqhiXMngfOX7pnfZ7zfy70RcADRUg7qP9UV/vo4NULc4Sx522/0
v0fbEB9jRUytQ/wgzdjTyGhhFGgTqo/n2VNjYpdV/kIBOrNK07Jseki9JBC486MshZ/5oNGmksLz
be14rxmKz+ugmJGNe67zRkMyQPzARXJL1BocW59N635NM3lioVqBr9TG9diEvqAbz5UqTGaPBWu8
1F2jeP72cuSbRxjpZqwzfvXpvSDSiY68cjbZ6WhZtXYLW1aVq/AP4TjpLekMoCrg7GDNeja8CH9M
tG38wOXolfik1m0A0KWOJ5VwcWQIknNO7w/BoCHcBfBCNPoJ7oxv5iXaFQrYvEXgcz5tC5iGXiWf
0NUP44e68ccJtzoH/k2N/CoxymQDztx/m5/Y41bgWnVPdW8Ze39E8U1W1CSs59pJyOXWx5JQhxo4
jkgR2k1K26Uu5xCkGTRgxvy43calAiS4Lay+IpcfyP20uloEk6lj4Jkeo8Ifa5PHKXHWFcQCHEqx
PMJ3+m9OUMXysDly9nvI5l9LnCEPzeixHRhTHEKY0o2nyucbKylBLioDZfEBfAOLP0uapZBP6OZ5
RYkhTILBrDFKKNF2E3mT7IW5ikgjIWltYnTNB90SJGnkGIaq/JOpLX5yBESUcWC/mgBgC7I9wX7f
KJSL6FlDh43lq/BBFRcWaq3K3tTQ0cC7Do3CbLg+A2txeuXKXWn0AY4pawUgHw2UX9fkb8VtxDp0
wttTymB9q+LsTLnqyv7PrnGtbniKsJS9/LdXYLanW7TQFjMNI+Lqto6lGX6DL1B1hdV1hMa0XXb7
/Iwkq4m0NDlAoV0p7W2KfZ5pEkjalMAJRZb0PolXazS+9K+W/WyL2kn97qQcbifv0J6HQT6C+Vgo
DWf4RuDnsJ+BGNgRbeVwAGbIhoTu4EIKDcR2z3eL67QbJw4bJj159gOX6HpOVKX6iAd8/xU+WIEW
TnJZJ3QUdHZKQGTE39Em8t3/gLuE6PqwYycRBsTH+e0SPz+HDgnT2RiZsRRKOe4XV9EeFkjhjbF/
zW5/0tIic9LSesZQrwgb9oxvfx3XO2CHoI0KjUvH8leRaTUx24n39qiJtxi+JAeIqyORbUM7K8Wa
FIQlIGu3Gp24aEAaTXAu7EgpYJ7uJ5XONk78t0iWdFXHaLkUvFgybKRFp5AEWDURkVgL9EO0bhxa
1cnLgDOlp9RGhInVYXBqaB3S0F91u4uJo7fnWcWavtYVchT36iEPRlQ5YtmYlSVe5prZELsTttST
JdeIYwh07iP+mHUngjp4Z/vxWMZFwGSBfYFG2XW18KGvqJt4UBeZnirh5+K8NPQwsm1KbZj43KGg
7Ql3yaWhXfZeRyExgQwUhx7C2QDRWKV78ySwsZhnqWOiMvagM6ak6sX6/FNfxXR6yOWd3PKLveTT
VI8MHSvM8PMUAR5nzZ2oWBB+fPRPL4YNH+KNsEBqnb0hwRUeYvz34v2VlhhkQv7qmLtfWQRU41eY
/qYZLi0HrHMYoapxOo68EOgo/6wxZnJdIjTIkXbr/7WDmgC53ygvZTPdJzRJEMLyocjeaznabqnO
44EvoTN85oWPw05SdE5JhMSa2UNXGvBmZ+mjtCPy23yMKvvgwX1UpV/ply/V980LdS0FDdyxOoZu
NPZnUWwoNyeiOoxtKNAKGZpQo7HCe60WCgzei+h99SF2qEYpOCHJLUnuLosEc2zu3vBjmnbTMNV4
P4qtfpttsykWrejw+vtCpJu9XIMoB65C8fiOGdRuO1V1gD6XI8wnoJFneCmXRpIIFU+NH1kqqrsd
CMiHPnDWzm0khyMrTZrCl5+KPqkK7nn8ByRi3iYNSdu5+vr6octLFPbcdlOgPG6PQxJ/V1GK6kyQ
Po5Wsr4P7eZQXeG0NDKZRTeAsQw1N1urQ+5U6rmYqNkyTUfiBQezM0EIR2j2CwAiOLesVK+Sx9GN
M8RrGG2aF1Np6J6JpGYlw1B7PRiCDeimYhKhfnYsB/nH/lVdgrjXnoAzK7J5RIyUR7FbqiwQ0GdX
wWtNJ2z1+csf4uog6kaslB5aFv8RETvGFMPO8zn67vb7d+msT8BOwnUoFQiN/zKVN+lO7mE370nr
aejs7nYpPoSJb7P75lblRrJVsmpCwVGX/onv1NbfYP/mvXY3RzFITAJSdpxlM+DPmUYX6KxGCRG0
D5c3ENdTomG+K7orhUxGHLY7Ek9y+1YtzF5pQ32Axl43eyZ5Zte9eUImCCQStHhORWTQwgELRtTb
0BTd6/VmeZUNOdqNwktB7gwKCvA2CF07EWSj1rOzL5Q25Qfq0s1/9+n4iJzvGJxkJwiSPI3zJL3D
CS8bZtBB1rDP+RVqF3GHpbnl6wORRYAVt0a7ZOvn07/wvyjoaRLPY/96NjS/QaEdgsrC+PgQ/ERq
EBmyHG5/Fq2R3YEFp7evyzlKwOBwgSjoS0Lbz+9zMBKWq5wl5o+sS0qKXkBr8kSmcx1bHaNtTE68
TXMUx5PCiHpB69NI4wePjk3bBaF+sSAbxQdm6ttMCyAziJKKGxMryRCxD0mcJ8n9EUWUxNZzVxcp
RIqg23cc3GkXVgQkdJNAOi9D1J7UQBDRpsp/LmPvkAlno/T6tv1OQLCj9Z1bkZfbN2xKJXKTmqWG
SA/Mn5ftYkPOBTW3TP2RBWUcIOTdmYW0N/qg/z76UXADPeoI78bBjDdMBgjdY8dB+IvUYQc84Qtm
DDR7JCHFSaVHYMULb8IewfyZ8X2eiQDgwiB6MaIVm6utrEEBqtNby4ufWX5LSfyS4FLFNmqgih4/
wkq+5Z7yBFdc3+GjqmRIuBcDyZSpDwHewZPTMSBMTp9j8tifHOF8Fbj9cS/JkQAPOxZ8AkhpWZJ1
BjDYcGiRqh84qFsn2VWkF078qxNDMylfJB/Pumilc5Kgd8zoplIWXKBWCy3uLb8G9QjWdlx69Pcj
45cdIoW7d7z4OIucNjbPqTdAj0rJrXCprWZMSz7hOpC3Rbbg93SXBhVVLr1Iry8p5OVt7UU3+Ygx
+yoM0Esa094V/albpBcLfvOIoGxz4l4MIPenfmplnOuh8GKoeUGOpemngkam+X9BTVEjd5hWpnsH
Nz9ySrPKFgw0EmnyddPQL+XdSRYqckiA5f4Qh+fY4wLbYQRlRLtYh0c0yLWXFQmcCF75RbA/ebRk
hTRQ8FIsu1EFNU4vpnmryZr/FUdSUvxQBv5AYo182QmXm0BhgdhIHX/g1Y2CjUn78wBQ5Dd5j0mC
GVDUEQRFKygVc8mmI17PvZuN7lWHC3gVBzynEovPRP/3uh1CMJaeSYI4R6zLJWVD7p14Oguw4fBm
rJjgKGWp6TXubVv4fh3kvK5DQb8RSUvWyuq66P8kmmqIxfIzTP6/fAkRC2aGbPdt9OP1Ozv2Gt9R
ODcg9GbYoEffiKLEm5/GQEwHItzgHASNlaU9npLJYlU0foTPaS0+E68U4hRUd572//6ehBME/JTe
HWkEWSRcz2y99TXCAewyzgFQbER0oeHVKHLkVfcKeTOLOxMU2Yqh7WZogB/vDeBRlFT0PHI+x3m0
l/W0LB8eTkFZsRZ7xYQohXYrhD78O+/P83DrM413nIxerkVCeBJ13E1+d0ztqRoMjHKP6myGfLJr
qHw5Z3l7AZyreq6vTxNCjsJRQ/TKFbjXdHbhQGxR1arlGghm4qxrR1T3gVwcFIuLyz4voQWWFaNz
EBMX9i1LbIhl4fXhDiZxx+gYy5Z9bTw3EsmiR0Rq/h02KDJbqltSHtdTkBbiainEjiUx3kuNjYR2
ajUdgNy01ikA3uGTIYwjtCpXwptaCC09AxKXUnmm1PpNHVaaBgJNUGrY07NrUpSg5kqIbmiQG5/a
9ZwCvxM8P/XZ/WuGMeqlNrei4Qi+2CBg0IUKnrzNG+F8dQ40k3Y1BbRQVlPjBJedQDLe/w/Ychz7
9jti1DOFma/ENb8wCMfTqsjlybkwD9AvD3AzO5/Tu7jpG7cLvjzGfsAE05A2Tazp0+sWJeqXhnw0
S7p5bme9uKjfxYHfdvw/lDEIBXqZVtwXUZdmh5bPjyysjqZk+ZF3hPwqpUL1HrhopiMk8GmG4xFs
M/g1PcLqDFzCbaYpk06T7dfW11NK/XS/blgBy2IxOX0TKa0Z1qZh7p5Agc/hP1S47ChvDtx2tAQc
6ht7sPY3BTrA8sh7nwy7eCjsBbri2JxXvJE5hWkBO3/frgbkSRpBZIjFs+KLtTXguRA5m6wqrX4C
F7rAerFpal1lJm/9bvGkSfsw3FGrhbLYsowDUGFznqktYHnNDbS4w8IW1IEtrfFpdrNc53SqSu2T
X7L7PSLlb/JvrbZJ0FNcUhQ+0w5jpYebIEZQyWvYltld+ywwMZjU2QqID411UbJvZyrUeeuJvqsJ
pWR5s9nKrdCQFSaecHSxCt6pClvtCn4jmE2Lcg0rSyhtA7k6hz9UFC6ecQgLfLXIFGSJFhOrEvef
MQFxaQaUKSMpAiaS28Zd5TWNtgHVejjv08axlNHP5o07XC/6Iu5y9LnGn5pd8YcFuUd81sVR7Tyl
IcrJqFMQxKynEikxGrPGCWmRta/vVFYnj4l2vkFYGmqzh9BjOaX570Lb7TMIEKaNNZkBYiC78G9M
PJqTc30Qvf+wvMVjPhfaAQvocqiFQmiQyo8tN8lCnX3l+PLxOr2h3JYzRVrZijn7LuODmgPm81gb
jsUIJhma0IMBkHxHMZekOXTDbQFoVJk6xHl8UHBtSspOLQdsJ4CzyQuGuzEI4NwUPpWXr6rxljTs
C4NWzoDekj6YWy2KBvZHY1FOIQDjdQmHuHmFbqzHyiByddkxaOrJPBENHuVkBE4719Q1Nyzzeprf
NvHbQFl7aOvGveKvCZSIHQlr708FwtWFGtuSuQMEiBnka6J5T3LyvzRjShkPwrtD2wq3RynaIHk3
o2hZEMDwwNt0xsUrbSk1sRx231UQqrcasoLxsyKHGBxoYRylTs21UW2MIl/j/8vC3VATeuqnUaGE
Se+r68tfmRxCInj38TMnNPjv44oi9wTCHRHTQ30lmwRNlMMcHlEOcExMIE6NYvrbmO/nr4UC7T7L
YCudr5Zi4nn8vQENRzNQrJ62+2ItkspBITz9KZz5d3qW2mebpSybPZxffeCz9B7POvUib+XGZMZq
qeVfqd7Mfrp17+rdj2hrz7dpeT2od3L2otJvrEXFVzGFLl/ZWS/g9iplyBV/UJ/esD84S+aUBT/9
U2ekGPCVFb9+f+mgqTwZOIChPH+c+kPB5eJJaO8AHx9iopHTT6putY6mW39l3TzZlgR9cydVU0zp
a0L0wh+tJd3HULuVP0wS+KawkS/mMyruwCJ3LxwZ/tkyFegW/zQdSn4dwx4jVOEIerpM5Sar7snF
1Bj6P3Odm1KF3FwilzsGcY7o6yloL2KYMehgNSnz0QwsvwgEAHVSySXLmM7BuMfrKd+i7MU6X3H2
9JrjpJrw0eZ5vNvdpo4Z2te3D7UXULNL1ms65vjFiRjEMUErQjKHRXPw4fYTvTgpWbKxl7Q+i2LN
hYIVFteEBV1uFD+kD1tQG+057lrSunLM3Kq9zdTCB3Kq0Yuo656KFXCdnkAhAdlBMbhU/UZWRUjN
Jki5kyDNMuAiGyaVr4AyTGwfI+aa2+8FypRsfUm7Aa6o89ZQJEBvwVk2Qtj65GTpN+G/vjSQy25G
rNqGCQujfx5i5MziVjSKVO+Wr/N8qNI/JkPDJy7Q/4nJu5uDlbP+jrfnMsgK5RTziyBK4TGFlbZX
FwOTF5hJviTKlwiB4PaIJG+CsHSilF5xhgPWHpVijDQ3qpsMhWR4eIkXN1qoYMXDFyMCC4h5vjBV
QTDjhCD6k3DALuQ07bygdJILdRO2p4knys2VcEpRjoi2XSPNm13O32AlvtJz1tu3295fkWkj8qlZ
lCUAfTFMiQfAOdQr3+NyttWy53kkmOBgjDFLuNMKjhhc9L2vLFtM9Tlh/6WPyeO4YVt4o60LGv9p
bE5AqLsVjaRNLxKGfM6wdErepTsLK9OuKrCBYvvJCI18c+vfFWnPWo9cSQ/o3ccGEhzXIHkjz0JV
ZxOSWyMOQDfr3ZrD6JvrjEfElVrN7Vg5sDtFVbotWi7TFiQxicVY5kVEMEsgdJ9nRBr/7P/jKCxh
4fVfZUU6+eN6Cr6NxGoOmEpxu/hqwaS8uVtd2pwW2U/ClFqwlPDHr+3EM1FGpHKb62dDdZ2iNej9
vYkHkP/CtbSFdRTUXLayWZx4zJkiN/WQxvCbLMfiFNsVNubgYE2MrwWVbCevjHezjLVanVlQRXck
834nkJ11jKbjVPyMCHLwE4LE1Y94KOMz6iqJGtXnm695V0UdnCf1LR7lnCErIedqGe3PmDYtpH0s
8uqD8eT4tzbmlCaLIcv67lPedo9PzCUvjz8SV1TgNvckS/4kphqvD3lU0WFq9Nsw2a7fnq7F+9OX
3CMtmnEUi07W+RJ4CMdgZUQqWGPktkqOT5seh8NycVH0AzOPGUfDvctz9YMu7kKlwpAV6Eq92TCs
0Cqd9oJfiu+i3laWGv9Yc4xyg9PyLlqQh5qrC1xB3582Z1FxHDqc+SZRwr8AQBIW0z4SRfy7yeB6
IQco5EM4GvKNTP1tXGPtpre/k+M1E4e/feX25AQjA1ukPkH7o/P1tll088g8fPL6+xe6BkUPmpET
l65pr17Iv1tMPQMkRLOVwDKCPwo/NF1pTbMvBzuGMStuLF8XYeIDdQaCl98r03/EtwxBjIMr5xkP
KK3rUMRE1rCenuS8dYSYovFNqnalNtiXpAFYV6c/N+Wzj1+6Fwz6ENOV7E9bb69SJoiXFCmv8LTh
78W6u8jKfFq9C+U0VVAOKbMqEI79EL09bDL1UU9ldh2k44JZyhe2209G/Ov7bO6omWrS2zwwhEpE
yJ/yGW8faEwuMOWvMQjN15hipnu9IIxMKAz6rpLfSdfPFrPt1hZ4+MlLXXDTJsxzEfGueO0ixO5h
mHjQH2AuWxJCKCaR0Fu41m3lD9Wc8E/bCRJJZaFBtZr6PXnjvaxIVyTdKJptot2Pfv4XBuJLkEbF
M61J7qBN55pWJeRDKbzMGtjpOhkm6m3VHSXeEhsJcuXGmDieFl4zPnIlqt+KT5XUJav/ySUpnSka
hYawV42fAWgq4Yae1jooPxrLK7LDwld5UOTkU6fC3J8EHmWXxGfqewxkIym4ivUN9600LB6Z0IlZ
MI77ExT7KkHXYaTSh8Z/DCqpIq7zxmhPSvsShB0L5AfTmc53iAG1JD0P3m80ycRP6X4SgCqhC3gQ
6yOSIokg5Iaw8JLntnZ6puxZ9ua8aMhorpb/azEighAi1WuNYoZ2L/eLLeeKQRkPsOWx4c+ZmSM3
ZUK43j3jiAw97vML7zK6tmW946QKyy4Rnqfor9V1OcXrZJQmfxFPKAwJ2rXFAbMdJaJWD9Zfh+iQ
pnh2xj2OuCQIuCDfajtkRjwuOol1OpLRSo/AAt/f773so52Q3kTs4TTNtu7wBaKF0Sw9UtiuQneo
++kXzrNICqSX+G1fwbAyPOVlaeJ/teESZ4rUfpXlzbKgM73jPValpBo4ni+rWSFKY2tRX7LHIrzB
59WfFOjvgpTGmLjtX3Y4UgalBamCg2MTujdUSmnYhSaz60SaL28EeUdhBVbYaW1jOhJuq+skHiUu
7y+S889Uqp3UQBE6ZR+5FhFjhb8oKh25xwgZARBpu9udkKiWHoGMI5z9duNV2Qkx8U/exwgYAujy
JtyUdFSQB/nQ1/GFVUJoYVkKkGelXstqUOf//pz+/SNxnCF7l3d1BIkG2TLaXRYyiTPysycvaMfj
+eAhooRaXE4YUsAhf0wFDG1B8iH1QEMkZUANTHmzKJMAIu9XzHNUUExeI9JiefF9/HBrnzTLUWgQ
N5cBL1j3OCifMhpFbXUxgieFjbFb0NoOQqY1vEnB4zWEOpboscZcR1EnVh0Mm26oao12uKi2HwjV
aPjyfLFZgid98qBM8kmsAn5kDdyuFStzfcmtzdoDPGKLM3hLqSjre9vrXz7sQSJOVbD24FiVHeo4
qP7dYQ7eBD863J6UAc2WYk2X+nAhmxguZdr7NO6l7xFeB8jJFlqcJc2xjAciCmu6rLhhrsJS3Vu1
/9SUA9nz7q3dQEgF5zVOKRpEUg38Cl/9QHK7EjP/aRih2tjPiJP/po0UpRgKfuR/iaW3iV7KSY6f
D+0fVg/fZ+118+PonVed06Fg6Jj4SqYldRXqEM4rIwwzO6DJncwbbswug+O3ZpnlIVrGaeAsB1od
OVxA+3Ae33rjV2iI7Vvs03SfRvhR+4ET8zkoyHu1byQyXTkXWkFf3LcXIZ6gDCeJ6eEQT/B9h3lY
M5i29OG0sY4ZtlY6AJcVSpdRKpu6twqsZLfKTCJWkfxX9wg3YIw2qsNpm3f32vyBtKUmpsQ0NzR1
yUGZf05K1UPGGCmf0uens6OBh5YH3TbPvSFh/mGbIbqLL/wBqOJhz7PUmupHVg0J5we7EDYr/sEt
Fp8KWClCblag54Jf+cIHvjwQ4YAI/ecE2XCWwtU8aOwAfb9M8Ul9nG4q8OKvO/O5BRs9BPY3bIOH
dQYW0Atk9v+yhBJ7XqUDCqmfHvi47ji2Lm7l2LJ6o/bMnkln7+zEVx1kpNSG1g1oYZT3TKdztrTq
N2F5RE7GfoJhLI+TCyYICS3NwPKp3wCR2zxNUbP6AOzTGEt4lDL5q4pbbUZ0t1Ij4fR77ZnbQ0PX
QWU1oUYfIBgO97An0zLeMc/q0snnw345X5LYkmxNw11ufARou4p9fmv0g4Na7ds/P+hWFCRHFjE5
ILp9SXWBO/fWuEQ37xD+gYa8wP/Y/7t33N50AhQWqVZtquFm5plSep+FWUkMfUfja/kaAxhy/IE1
V5r6TaTKaNa3lcMz5PdsYKgm/asoSS7/r1n9gmmD7yYqTGu4/rVUeVQjilm77Jbe6Q92bsFtRTW6
bBouBbGWfJ5Mc859Kg2IaKdYjuup5046JB0VjbD86MIHxsUOJlSmk5/ylt+Xx+y4UmL5PUoK0dJR
z1Y5SCNGH77gAsHJVdJ1/0aOA30KXOIcKHaymcdCD8qYUJBC+9UCs7DLbObaXEIQHbbnoVUpI5P1
5jETqW2Fqr/0sPuQ+cHr2GlwnteHO9LPBuOgvgMUEYqn5uIaTBB3zeeAq+zdMnBExw7kQRQmbkY7
V4syJ/dhYRKpFY67ABFsjavHB6W40Ew3FdSIMaMUDfmFVjDpDrDX48leUeNRlhaTSjHcv2BpEydq
7eK2DT5qCPjpHxbKvVE6xE8shbKiy6iFNvlAOQ3M1wq/Z24CM36DErqdFAVX69iYOkzuVoIj3gCZ
/Kelh6UeYfv92HPwo0R2302dJ8dkXx7RESdk2a4ei4TJqPAbCHvio8yuKStyijMT7p7m7L1Ro/+6
V+oV5MjTi5PwVYEvh05QPO4rO23JrC95W0FCRaXsrMRKeEbflH9yIqvbdJEaJp9dP3Vb/vMlHnOW
3PDwpFv0cqEYpQUfEnnxuCUaLh3QfND6frOjM+MNrT+qp0NdZ/RhRipckYkne5PG99tLYb3ptyvW
A4CIWcfKH0Lfac26JwtCU7+dPvdTXKYPmdaZpBERTOaJJcXAZzdC8ShRVfyGznE1n/nyaYR6PfqJ
2qvA//HoWze7G+8KvG3iI9HS0u1AKYo5z9GZtwMcMLQe0QtJStIUWUlKU+DuI4s+PJ8ue/tiOtlL
3w5jNQqyiaLNkjVm/Lt/dqq3l5bqpk/b6CDJXp+YpW+HZpxRJhVW5mJFVNL2+SQfAjgSX0XzX1Sb
iB9Sr6QJNVuEuNPjyohxaMp4CiW+UplMSxajvUAWT2s/igZ4dS0DYwZEoE/qBZyTykFOeuIWlH02
vnRBlRi7gS+DQFri21vjoEz+Uj2uzyZ/5pYMl4QynKraGk/vKI3mybJZFiRk+2a+sg0K9daLegPz
OBzTKZczjC+N6Lem9hxrfuKvh3e53gyq6t705RGzJ/R1rKBOLXVmKg981Ueri7vPc3TZodOYnGl6
vdpLcocfgDKZcCy1DvqIuwebKEEdGYPB969xTfdqVF30zWUYE2BJBq3CLrz/4mGwPS91T1m/qYEX
InABgXUQqDd9LxQOHV3gy98yZwTGPf7HKK265KjUk8ELkQKqwZpwiIdjimAbcW50sSVObMR2OECM
jRi3sUt2HoMsE6JSrHTFfHnrm2wSw3mu6NlAnbrw+odfyJoBPWXip7h1+ZTjmBDUCL81ZjLh4wp/
pPweLZEnIlF825764mOiBwAM5r33YjmLmQggbprbmSRuw816NsaQ3okoZ1Bzl+VZsjYeCRV+jFI/
AXZtFVJ1Q2JqC6WtFxnVJSkl4fVHHI9l6wrqM5cLXL3bf6o/sj5IaHobbYw6zLVXjgkBg6Y7Am0B
p7caKS1W9JRxDBLd9gjKF7mntGbvR7MAF4jkj3iKytyslx0h73JGQy/mPV9Popv09Dg5IX2WEzNO
16uqAfZrDLInQskz8LlH4EVGEWIVKN2bGF7LudyefHE/+KR/q2+emlNXKRw3OwQfouf8YGDh4x/l
BxQ/+8ZgrGvHo1cLOeRggX4p7Djz6BZRmsAMeOk4RchUOTtzRluoJ8lEsE3z558oHvYP1RvPEaBH
9ysPFi2Vt1cy6+DUqmDFD8wBvfq4rwxnqoQ5ZVu3ZFXF09Mbdphc5pTyNzGj4hb4e9Y4kc6CTohV
FdnXIwKDpIXXukqlAjgKf7ibpv+LAFX1iE1kfbDa1To+TS1r2MvY2mYYXG1jRpL7pVvF1nhxj6qy
k+Rur9ktdSKjSKCwm2IkcA6K4yYmn78MDBMV6gF952Efh5QUahEbp76D1yqQUQN/oaQPC1h6u9vW
eRHm2LiD1On5y4bVTJ1v0jSfQlhDlz3IfT2j/FTaU2plXJ8NetS4C9InNeS4o3y/tYVjQ8L2xptK
FX5BCZSsQxCaVrWqR3Kj7gc0gK0I9QkHqBnFdpRBgUgyiZ9PmkH4QvfK4QhdHQT6CiJoHzZrdYzK
78qIo8xUqMyntz/o/VJdpA4Ffpa6KIzSUx/VXXUXAcLEOT4Sy52MHXJmroHJNSVItPsqMUS6En6v
46vONr4bDCr1iGMyPWyLaP7bGo3VgxBCSNs2IQ4v1a9MNNb6i5vzG8saYkg1ZirGYhp3Trq8DahD
0jfkPRb6cH8gOv1wWGNTxq+JksUxFQz32zoRy+ClBnznIyVmHOT+c+m8MAq1tAzdoxMtRKODAQEE
MSaKg1lK4PJCqaExR6dJoqoQFfwXktgcGPQAQkroT+hs2c6cThnNQtvtr8/tMqP5N3rY1yj5oU91
TU/prDsLYVJ6pm2MyOe6WPQ1LVFz5lSZyMnGpQS0yJi8D1oRS89vcnSrZDdWcZcAiFPmuCSV7NDg
BTyjnsXEPdNjhFLr7gmSuIQyNSWRX9x1LAoKU8iKivl/sDbspRBQ8IBRJ9wFUlyS2oXGN2pRs2Ml
xSvYI3HGS9RuZzzPrDoEn5YbyqJOA25EkJwdVSMetoIHb8BjO13TOTeePM+Z3U0WXVi+CicYaG9h
ikUCLe9yz0TQvkme8PvETwYVxsnSxzQoKmjLr8Plts+eYUme5gLwkRJX9dWMZvxjKqXxMzdqoYTt
gQMLIiNym4Aobrur9mDcgMadvxpSH4LN/9LE0ZIs+BFkk+DyNW2vIeJJkTgvGtVDlNSJIfgxW8cu
QAfwUBvvwIebZed0yO3RdI30iIVxx+PD9+qOoSRMWPz3JbAyxSoD0NbNCE+NFJAWMV1Ztx9BqoPB
R3aIxSIYPF6CUmIl1FqIeOCJKjKz6KdXj4GVJIEigMbsC4oM/IzSQ9rRH5x7mIvK22EnhNopSuLF
Bhsf1c42SfmrCmzk/0aedk+CIoxraDvzAA/ahJzC1oD3Iq0thT4Px1uTG8tbupzgUZGbuTYeN5c5
UmE2uh3z/SZBbTU7K4ju0faWp4is92BUeh7PwRrIKlf25V7n9OmHuT8oHuCqDcIM94T0d0inkfCo
ogN64Ekmq+8X+PEuT+FzCFyi79URUjMpre7n9j2Otcnxfnb/jWTaWhy44+nunf8AdidEPDDwO2qh
ZqZWf7MAnN86c1Zcu2FtbX0UxNhdWTiZ9EFwtxEiBijKO9hrseo5SjxusTRrvpmmr8BJF57oDHkF
a9IpN/XNOzBXY41+62/4l0m+XGWDciuny3KPP3Bmkkmq4rv6WSaZKi1c9so3NbiGskD58Jg8wgRN
AV6QDAwXHGWQZ/LDzDpW3adOkchbU2GdmcxxPtozXmozpE0YrArQtVjHJjAV4Oy4HipXPuSytMeP
JDQE6lJ+AkWx4h9/epW1O2cTCDmrfGNpx3ayW3AVBdnhp8fqKFX1Tw4+Go76dRdNJ0c8egCSpGME
SK02Qiv/m/HSbSW3cVv8h2PHAUXkA7bir3rE8dfBkOjWO45ui/rYJ/0/0gzltSIuEVgy7UD1JW08
7t12u2H/QCitNUXlYxWMT4wLAKPQ5kldb27IyePXviXPaEJmIgdwXVkv9XLul0HF/Z2EYcHNgYRV
CzT1p/RoA8HFA+OJ/z94PYa31bUx8tjYr1W0rTEHYlsDgu82u9/gs8KfsDVFnR7powvsh8fKwKBa
sE2KYvMa5rd3hPNAKakMWtldhGwqXPJKQPTd8OM6KC5wOnw9u7y5dB/ZvzZcvgOfbuLj+NHapSnI
woVtqzKHNO7xcNOoj/ddcP9v780Wp/WlUDHHGoG74HGvDomcyDxPLuMt+h3RKLVylmBDUV4OMG3d
abzwJEOAZP8bV3WsmhnVhs1Iue/Pw+qFqi9MXIXeOmztKLdQEOkZAkcndCCUibDYzOHpS98psuD0
3rY0PPjGK85OuJWUHHVzv6mR0SQBNrAj1xthEo8Jc+hiH9abBv+73BaiLf/l8wVAqYh4hqxTih4P
SMNwsc6dfOLvJOLBRschrmWDIbv44TDBUf5QbWkZaYB+9U35PqP/rX8U2u4qN2UePBF/czbiAaGA
RuBSbV6a3Ej+E1LEgdtoRlVdHmS39E6tkxJ31LOnw0G1QazWlJ3R/3XyALy25ogNFwyOpCZuLYPc
BfJsNr2P/HOQXnp29DZEsG9Dgf2Y3qOZR2MMsbiS7r+3ZJc0e5iQq7Ux6gsAs0w+w7Lw2btEftP7
SSyUYsFMTnbSAInsuOXJb8yzgc4pWh4frmQfd157xL5g6Ne14jtX9gsSufE5ocXeFMJXh5TIk1fO
3ZJo+vnItVslVVdJ6JvIiKn8EVA/uWUc45xE8rhFpTRljmZQuEjZdF1zrBC5tSzm0RJY19Bt+byR
68jl1gnMpMgV8T5+LbREP1N9kj0Qr+i6O8Pbiv7w5uvg0POuNxgm3ABhrCmRuOHT/yCsnnvOI+fN
qx0zlkwumQvyAfLXNumZrUKv1Wh9kEOzrjrB0+UeCbCrLQNswtEknHz5Qg4wh9vyU/vQvoI5/61K
RqaCRq1sux5ithlNZlvxFWJJCZZO8587NQ1exp5RKhQvaTd3eAqAh/G7KAbp4ZuAWvnFspNwYh/4
nyIGThDfkq+6KcQa+uEg8rz17oI8nbiYHThISCDlHINOXetAC/54CdAKrHPFdyGeht1zaYHs0bli
r/A0j8Rtt80KoMxOXBygAXhv2H2E8Y5emxIUGN/hx5XzJtQ0boQiCsUV/iUdy2wKZJhI/gy9CKuH
F9qxvcpNUXe0m2mcnWWPTubfHuDv0G1StdMdIvhRXh7bT5I7uvd1rWB/OZ7w6S9tpORqSn7lKU4Q
d0EyMR/NH5gldYMg9pX/xaTywVy3SPYIs3KxZA051UYgwgGcOeAothpU1nMg5/kXwkQVGZEBQeOn
2MhtKcCHIjUKCW0yy9f9rVfDWKC21h8XgG0i2nyT4ZA02iyaDyW9rRsQegxlFMleErv3pHD8n54d
rEGe6jUPXH8Wmvdzxg0gmK1WBx3wZRXKVdH0kLcnPwQlxVIlXnE0PXTHKQk3Mmx4MuYfG/tYGaVk
nJU+9gCkwJv49aPunryUYwjglTbepW64ZSAHgeQVIxXlm9GMfZufkb9Xk5/OLE7B9qch8OuAhrZd
oweMUkF4DPKFgmYbg3xjlzcT27N2hszewdozLaWOqoS4XbKqlJkyE3eWpU+WQ5vK6aYTVL/JhTj+
m6ylxGuUFcwwl7MtoIMfm8M/UnpByuWCgZL7exVplEQHSZuNakJ2mtCKFjWZ5ZM2qTckuowBJT9f
Vu6DZxvgUEoX58RLFt7AL62kJtXsLHz7ONWt8Y6VNjYAtgTVcCfMa+xj7xm4nHgwYaSe0YlNydEK
hNb5VoTMzx/xzj/QygjTpBxPGxIAEHCtqLiCsg8s1m3Vel1fidp6IcE6Hz2yCd6Xw/C7rL7l1z8d
orFRaXBBtOqtVMNvBEPzcGkNR1XDPg/1HhGAb4fy5AY8NUhY8ZAz8m0ithO0BF0ws3eQkVaQnmb6
XmwZSb3jOyfUmXJoZJuj8tyaqMpjIrzgWTfrgDmFx2p++QesM+X4X6fPrAUWMevYVUxFa/GqjNkm
AcBVH7ylJ5O4eZVzwenNtLnXerCTauaH3CBiTC4205N6e5KCRrQzB7FKG6fvHDIDJmdabg+LkVWI
oO06+ld/f3LE8NDtzlXkH6T6+rMnENhDmhy8hwT3SHBtt/OKjvAiGF2603GRyqjNU4UXVG66wjXJ
pVaOF9TOi58ZRqjra8W45jNzKoVwVBy9uEG5dhA7XdGluYhL7d0bmz6LuAMi+xotmt7WZfs7X3um
XFpvWAl+EyoNoCD4w+ue4jkjiaIS0nLcqTvebnGra2hTYJxQedrrF85vceZ+KCopytCXlr5BAb3n
pNC5Im1zgdwP8H9kKMH4SPGgmbxzs7RVD7Uk6N6bu+5S6lVNrM86T9hVIaiY76XR8P+t/k6u3DJa
elXgC5dDfAY6BFHsfVjNqtzoTr66b8Ad8c/rwKalKRFvgsUU4nw8XmUGOJxNHffgqT5GecaK/0bK
ixi1FCYL3/+YjAJ0h47j0HqgV0P9G3bi81wPYWqvkKPzQcZ8y2pDVbjoVpeP/HtBnP1MCq6S9X4o
2l4Fgiq+nCLlQWjRS+55Ykl6B9d6H8OXaZScXSnspQCXjjaxvF5ZMClMaAG97lYPIZJqJ9SB4yiY
nnqg575WGBG9GFBA8gbMZ4Z0yXxXX0DTQYqFl4KGSJiaeEkbdXxI5Z8p2e2N/W5uIMNOYd5ob67q
miSlixPcUeVW1Uew38tVSCN1D3JNST67ZZDM2wRxmDhUOF7+Jm5oPH+cm7NEPbVbAWk/qj5p4enW
Y2YLniGoj0y2d5IFS+TX4k+AS1q87oXTBI1IgltdxDopBluwUOy4mMsNFExEwm/SEcinDpdfM6IS
7DjEzPfmXEtRWwBfDFefWwbn6xC9aco0Swr7hPmpo+j3LaR6yP8c2e9RPF7ApFBj3b9FVlnHapNi
T5fx1GZZQN/msm4Dg7htGzLm6y1KwYS8eYeEcr7Veec23Vcf9SchdWMMAaR1DYHEt8iXhzHV5ccH
nyrpHQpXJM8/Pl32dDJ+je7BiVeh9APFFZDwOE1PgUUTeY5Gd9G1yPIout8SzM2PEnHy0+DIsWDr
a5VfHGyPLegq2WU7iL1Xc1lTvI+Oe0fZtF+KF67GZ8WsBWlqecM128ps56+F9kIxMVfNuzdflJmB
aRj5eIxaQL7VoK9IpFRnNgcqLnyMQGsiO71KtcoVClOsvZ474FF/183J1WSL7zC5oeqLa+0u1KfE
zdFQFQD/m6N2R4yv9006uGU5pExCXHdpUmPCP5zeYDnUIW2cw0ovD3CzbX8lImcMKH2pAWI0c2Jn
OtxpYve7/0yPN0pPchlMz3QVbRWqRTd7ynEQTFbk4/DUW1CB6yDBt1b3rFupZyxXTzqOeH3dTfiG
0EDOWVuc0PQ7nMxy1z4fOyiM7rnuiSdC9a0rpKPi+u6Ow60QR1Vge8CXn2YgjQV0qEgVReIQkaW9
dI5QP0Lp7SB9v9QuIh3LZ268Vz1OOankViwrW5bn0aak4uygRWDoOiDjajaitq3qwJTphcQ7GUlC
K/fbx31ZXQeaR3aQHEV3n5pLLb9rLg+INkpGlvjDOplUgDq/+EEXCq7CenowjnhQtDxxgVRiDpgc
jYNf+V2NLXeYqQBi27aOfoEbasljBtVK6k9gY1SkeXThEnzHDveFM6Njgaccskh9L++mhELRWGSR
NwNaJCVPcQKVNp/Ia2XwXsOesnbfma0RCkA5p7mNleoCL3iW0RcZLtrZ7sbAVfBJmtIQDGBxkXhO
E+CA6g4mqT7HSUcHZcFETfzrgaqSdpmx6qnjWFuTi01H8Pb4Uj/r3Kch0zjGzLYmch6rJnyf9TBY
ErDq5sW+am3ZzFeyWogsI/HPHsjd8LPwYFyvIdNdcYk63ccstcVWMstO07XVmWJObaPIxphHqXlu
irp5YWqksg6zzJXbbwhMPcLHOopbykE84rksqBSiUGFQGacEuVt+DwQ3jG+HerMzt5i1v2CZdKhI
qKCRuZKTBNb76gYtj2CRR4jtWwAOLhualv3jEvTD33GMCzlDHjE+v5E4LPjXo/hRl5+ebd5AigWw
0cKNnvYKDYRx/UXowXnQj0YNbTgnn8lxSu3QwZDiyqu3FGPgYyaxWlC4HZXXfu79vBd0x9LxBors
TwH47F9zASzzDrjTIM8UGMthRC32Jv2l3PwGb1DlAhfb+izC3wUfcxafzauFwZHxu3niQ9DMqbIc
RwXf9LV5exAZ5OCNukdJpd8skXvnVdMfaowDh5gI/DMC1U+N47Q8GbjHONJ9R163BbfYqxMbD+eL
wHklgACt1cs8G2zen31/1W6649xh5FkbGSheM5ozv3hYLumMfvAgjajv9TMRFP1rzdQ7OCwb0YPS
6ML5OJCYuvGx5s6d99NtzvhVDbst/+xyDLx+zcB1GdQinbYp4ZUwLeaFhVE2AAS3GsXTXzvbqtZt
wUCGERXCdQpC+Q8ufryxjNxuAYrMopYdJnkuKB5vNDAcRLOyvt/9lz5kszwKKyJ2SjLHJeqrsfL/
KtmdiY5VlaOrc0AWyI/upAWHk/EXj7epR9klrUZ9LjkD/0QOeKDdz+aKC3dcRgs0NHdPXtbWb7X9
YY/Rqd1FPDyquhb86yxJMBsYJ5+wzex+5XHd9TUCKEsU/OV9zYVPRMaT46F/evZUPZA560ZmhPNa
Z0h2bvYYzNLSVeX0zQw+yPQkkK1LZNdTOFJ9dqhj2GC2FWK+EvDOpam+BKp816zp53pfzZG+un9z
t09Ecn11dTRrvo56z9jevvCo0njMzVQtrVcDT866OZhCNt4f51KxU43EjlcwKKIferdn9s4FUhP8
9UKozrYimMh81hj+N51r9irha7yn0/1/SZJSEJJhnj01jBG70jUFfbT/CXe4EJBcaXB4Y4vuJELg
/j2q9MZ7Uuqifr4S8fIvwQANFXOcZKZWf9y0I6w/zppO31MGNw0CsJXgaVpPE62CIL5WjABOlakg
r47JW9GXlC60lWCXby+ofm3G7KVeT3Sh1QVcEUmAhlzhES5SvHv8oXN9EjutssF/B8oS9h50TTvv
F9UtCvGHRPDraZgpRc9Q4CE765pFk2KzmyvCwwBOBJ2VMdp+8HQMifaMQ9NqUnaqDbWBi5NHH8o0
xUNAt7alcYUmzHA0SLgrKmqjVdeSzvoy5OnCTuVg2DFD3WSr3T2yTuxTG6kZVgMt9+6GEujuqYHi
KTYaQisEd3s0bqWpos0cvzSFJNI7QV+rRoqFZhM+7dyf4B9cGlPdzoj+aaa+jg5PdyPbjLLxW6Zy
Erh2W7HK8NxbW6e+dnHjGAxLnDCBztfoNeL2Vk8h9jg8BMH5Hk+d40bU3KYAk0bnrBblAey0Xsor
IL9/ZiH6S0Obw5kkub76OC5vDXh/GXOFfMLS/RGIbNCk/BhTAtlvN7UX5VtfN7dtHo/36xh+Z0pj
/oc+H1jK2Jw9Ia7ADdQrb0U5zf1o45sIV2GT3ruoWGZhbEhgazJcXvhpHwrXZPqVpVwpv7otcyHc
dqfwDNXHCFryiGh/STxIhcPN6a/U6G5r2xdwWj2bS8d6t/dy3dgyWeLkNmKEhGQcY5G0FrWLrFm2
dAZXaPuu9gcaJ6Ad8/se7+AL8R7nF2bk/hsZkM7nTp3NEpgNq46MDfHtcuaRkvshVbCC1jkn4NjA
ZxiOIy+tVaqLkHIqy3Y6q8MfltBA0Y1eicyLCjcwoij9lWxq9lDKBcGr0b17EjlciIx6j7NqEOg5
le/9cY3lOZP8T/4yI6BLHsDKMLNZafNlHipx6CezCwYE1p48cRwAXccFKU/tPehXa74/akn7b0t4
qjiLJnmfWRP2BPwXJvJ2NiMST31a54n7A/sYJXQnUUMzfHZvbg41tS6HQespRSqo4hOZgJLq0FjY
4P4hEf/iG3O7KqBPki48hVBVPW1ZhXJ02O/9vZoTWEeDqfKA+E+bUt60gw26++/LKYdX4OXTbUDS
cLebKcDmWRAXFJteM+bzYgJdsU8pKa+dOkXWYETzCYPmz0+obmJxCdXDcA6NUBl/+4sOVbXDwlLo
b+phskHRvjtaEnZlIYIJUKnqSlH3VDTW1cK9uJfyQV7BLxZNDLF6K+zRZW+v2VoYQMJ0R2fWJiKs
8CJI9SARY5yccR7UG+wwVJI2hwvJbwuawExI2g4u8UVAWLLWXbjJeXmRXYgs5I5gR8x7O+2Ohw+U
EbTo4gmonLIXO0U8y4iOrQEgRJna9wAphlSnP8sMBEKB0ufskydq4uH0lKkZHAprcrFuQcO25e4N
mw6jRTVPArPRKHP3fLBpQZICEddqNnVN96ECinbwiv5nCRES/qMiJWQV1JV8VcZTCNdgWFufFxdg
IVxyIf+L1wCy2Zw6jqU091O/zPopdz4sL9yD3Dg09h2qU5JFFEePkmGyO3ZXf/Q31Rm9E6H/11Rg
RALy6C/O3/Gmzj248ndrmE/Dti1GC+sqJ6BVEiOF9SM/XABojw/EDNy67sCe31MiXlui6RL2llci
qls+MjROz/UMp+7EccV8GrnKsZTeOWKGYICixQyAyb4m/1vuyDToZpRTrRHWqjo/t3+DV4vWsMC9
Pmk+sMWfdkJJWtlLOHS4ZrimjTigdPdbDvoUfG0i2On1oSz6ltCOwYOISqL1BEwf4NuqSUXxeIWN
eSg46N3Hy6j/+H1jiS5NG0PoBL0/LT8RuuX2ynTja9djhPWs/dg/PPxpvgAlITFpyIR1tuS5AeNW
c08R8lVVcctKJ9q2GP2tJSUayO7bHbEibmu7YTMYOjwqGjW+6SCeSYjRIriaDxhB5KB8n4gJNHE1
dnE0EKvFADmGIaXiKfISd4BWbH3pIm36NpCn9cAaZD4fRvqRquINjLjAgyAo2oTRVgX1jI4Ho/i/
WmykfT9xp+rVqqeuI8XhBsBeFqHsLRFJb+3AEOzityobu2S2vH9DlSTlXPq9920h6FNnjlw2G6FD
zAlgqLxHDnUn02D/0YSdFOnG0ZJcuM4BTAAVroHzguuu9uc59DvhWpsP//6QxarYZlKlUvSes1os
ort6HcKMs7gdEQ2bp1cJ9f8Yhf2aiSK+hpgrNgHVz+m8vKXgM3zUbmhl3thmcwqVO9P388PY/tly
EHEKbItLr8mNuiLR+upijDgwwKVG/j35yK4DnfqZ7+pzXko3e+u8oU1wCk35HcVwig+zwe9Yfur6
v1FsurJjyIIF0oS9el0xU5qnV/+7YrXs7koQEN6YL9sOkRVMxjk3S1kGHT1JuP7ApnazDjL+8Owm
sJh6DuedoOQubX19eyD7BubK5xDWURUI/MIpTIbKmKRAa6IMI2z7zp8nkXMmsPy/QFtRw2jEtNlw
KO/exETcGjlrphdTAYu8wuMXWrZDQkaw56HpKgG2zSx+Y90mhVA9iBn6zH8omYtD91uSpoyyNnNj
NITRRximIJ5eh99tb3k5qXlTeKqDRtbrzwkc74eeZ3fFTvRY6sOihNKY6Wr0tW53TE4tK6QpijWR
FatFaSi0Tluq7EMn3S4GCOeH4MYeXRCUB0FyRPYammc9+Ot3OPyI9k6PkNOQ5gKSFSU1FKXAt0HJ
r0a50xYKzjjJUVJidy0X7eZmsZ8WXbzTC+6iPqvhrnLYnqieah/PGq4EsE1aZUTCofdwBGFCgU7H
XNYuUhIDgQlc4EMAfwBgWrztHdDik5Te0fJNKwv98k8FHf84530bfOB1NFNC0nuyBcy0EYRWJSGp
FXtt5/6DaAlydrQyXFJMgOOwfLUYhewCqn7c1L0EzGOrOZitHCpWRbTDM9yuffVxqkpVDxZ+ir0R
mdQWqlx8QevNQu1nzDcRiemEwxR1ZAxLZwViKfcThv1IOcGeF+oH9wjHR+hYYsNvBLU036tEJZ4H
ZNCRs6wHONpWpILzD6CuXX9dJIFfYCKOGYq1hNXv/qsmPMbjNmqrVPmtU93F2xsYVSuExI9jH5cC
+5fLYkuXIPfLMNlS4hRVhIplVZ1ZVJcZkCgRuEcJJL1qmvI44ImYUz9u43if+8fjM2rkM+Oes5Za
174ho1CdOLbi8lJY15XIWRNseWx5L8rIts6ANLX2k2Tg9ZB0sCWMT2CrqBoIyD/nKaRNiH41bnBG
XWJXFwGnU/jcXKXiRJHwg4vXGZVcYcN+i+oMpB1eE/cG8r/xqLbkiBeJIBP+Q4x1WcmDjivAlip0
vSlKrKtEjk+eizRXaTKaHq4u4p3sFMbsCw/iCdbsUTTwVuLCXrXwny8xGdES5rlk9te2EgWim7i5
22A1hpQgCBf6Kqvb4ZdoBtKQobM+giFuDglcEczh95oDiqLBGXmtntCvSwhLd0Ntbwx/eGcDbnrV
rrWBxUy0zqi8+CgCyDMgJ0+J5vkQ7sErGAbMpeXnkL8lvNDDCQc3kYbZJVeiPArzK3kgcPySAbEX
0e8zYwfwfI3rScIz0cwmC7eMbY8iLDVl+xeulf6AzBagI8QhTJ6t5y0P5rkxghfnOvBpBOZYBzjp
WU+lpPux5m2/k6pIafPaRKFZHyZr6+XQ7slBvmkZJkfmKXNIH89Mzn3d3qCvhIADycE6smZrl7Nk
Gc7Qq0pIQKfYL2TJ6xPqgJHUqYcLXUE8u+rRA0PpMjv7B1u8VRXzOD1hj7H6d3j9gO+4hmvGRJzf
wo0LMbjGM8B9RoDItdFNdyovfSPHQtuxSoXRV6UBIXQs/lHAfBL50T3rZDU/mYew9CwDb863K2UH
G2ubcLPOZCndimZi/oEhamCAjkiN5c4HA6BInz5+xHlR/TCzQE3JP738zBj5nao4HVmplFfOtPcr
lz7VL/swzgwII3PQZMg7EvAcq1qeVkub4UyXwlQa5kTjVDTOMtfgf62dLiyywmW+TZ+Yak0PqIUM
s8V7HrKdKR4mLi9dKBGpNCN4fKpB2FRB7GzylXxQg02Cb4QBYpSrGin9+LqzC8jI5jqS/HjLTVcf
Id05S2EdjbKSTznt+f+X/oCgNnY1i9bDiR+E7KaUyT8pk0680oIHC07/Kg2RU8zmczTsBJ6RHeSp
nFfDCV6IjGJhI0G50ScDpR27zSzn4ZQzVgZ6Yzk4m73NjhVjYw/GfnKxZBM2Bs3V6FyN4uUwTIkE
DLWUKeDNgM7haVWIB1kKhxooJ5QDQomJORndSPyGPhdLRYho4yjRIy+JCbFRKEmaVCHyHfgEIhBv
Cjy2ytd8Hp/odkaqMx5sfKt3P//1yrsZ4Zq5WATwNPS0QkFGcUAow559plsYVgnE0YB1mS/LnxpX
ij/JA7ElTzaGciJB8BdbGNnkaTmIW3GArCoJtAgo72Lif1/LK5JQtzlVylDcMs9/QAj816kzOWAn
lvhS7xJ647H8zwuk9TGZz7cNUVOG/zU8SC8nsw0ZvpR5UcqlsNKU+EN54SZawmuGSkutuM2S0nX6
+XUsQ7Uq2bNGEOZNPIBKRp7YqNDzFOKe9yITuFJVoHDna0Cz8IlXbIXMikT/mNAb43MvZrBOr9P8
w5rld2qj6ICCNz0w8XLKukjmIG0N0Ik+/+jFsS1Fr/PZAIcRp2OAHXRr80k+TFpVbPYiOAFuqRYl
u6ZkAmQY6m6zTSYqZtliOiWWd+rOJqdoqjWi6JENCa5Lx3Vx/aHzHvfiBgriWGve8rswCS2it3Nz
18lB/ZTmWWaQa1zvHkXHMI7hgcna1CxzkPF9QoMpzcpTcgFDoLEbK2Tgr9VBJX8Jn0uhTTa/zyxD
3nUMbYTikW78XSyE7mCMGpQjGM+UMTkSwB0tuNuvsJLB+12skf170vb3+NCy5SijlBbNiZddQ5yM
wb5n8QJCi7uEbd1vIWpkFMHHnrVZ+on00ycaTIxe7L5HXnYMmOx2CCRXSd8etxGPwqjN0xNg0SFN
JbDvfKvUFfh3trcJW2T2F2R5PghadMZAFlMUZ2Wv+Inxoe7P60i05OH4ZsMqD+utjk/rPp5oMcAa
0u4QUQ9Lf7Vbab1zF5/u4mWbQjPs+khUkWWyUojKxuULkDeFqnFFzxtDBkxAFBAyJ3T3QRmKPAnU
I8Q0AQGh1lk0/32pgP7AJElQDiJ/PDejuQb1t3oKFv81WATXwixZiTSc/IaDDM7l168UNf2BuECn
lFkbBjk4WhS1hjYhrPLrPWLkoYqX0yn9D8vYhJ9DpGHYpRQkjvUcaQcfAS75HVmV1ZyxG6C9tFlL
vaMdP8+zB1EIZDND0eULagtOpFHv3eaMtZDd51vrl2ilaQ1O7hXy2ddYXB+QO1IJOJNOVZ0KmnAG
UOITVvPqgi2rh4TymbU5/jQWVFYMaIf4Hq8tANRmU33b/ole4n8eNx3iumx7M2MrtDEzwT8g9MUL
ylaigs2U99+R3poXBx1y/k4lY5++gHrSQDo4YIZbKnPPb/c6us1g9tNdyiqVgW+0KN2VJ5C++5C8
6E4f7kMRibW0IKkVdYhJ63fENYF11+JtXOTw3IzMscqPa6c++7J9Br+e9LTB6igcehtjmveBNM8A
YZcAPLiJkpA8vSphWC8IU6NqO0R7ylocZn8DKhnB46LSlj75i6/R9PxLaVe89usbXaX46UaVDcYD
ocP+mtWarjI9gqTAqKB/MK/dD/DbkM4c9dsRQLsvM7srLrEifPa/DGCBdjVTMv1Qp8v2+rQSxf/O
cV0A1YTYPFNfjBSfAafE1aOZEPIQnboSeIYNjLaEYXmAAwHloD7X6WUyIQp2acGzi0vB6FlFohsV
fZQL2Jp77fBWnwCx/akpSJhrw2W8SujVFKw1gtGX9ggrWP9NmCS4531HcSniiGVdXsvKJ7tXQED2
WxHsWn5OKedq9MFi81po0YPjxCt+UbKXk8BUZTy4U8f7eWQqZg56VjpHtF9B5MmJWhgf9I29kY7p
BxJvojKtE7FMD/FJnG8+QWIXWe+YBDiVaYg3oVHSJR36zYZ423aFborKG8z4bsIu1IjzrvCFOcVJ
KCB6V9yL2gKLwEvZBojo4rpFuremQekZ1nqrFAUkiYlQLqjuY4dcngpJO8E2hUhaXhUmhlPs0YwG
OLdPlvGO3WP02aETZzjhWyyv1j0pXR7Sw6yBEwhr6BbmlcL+p+2aviksV05EUTmLHQ9mT9E+6mIq
K//OhlSamnB1s7IQn6woOpsyhLx3TVHOTE2zFJeI5NW15dJRI4r5oQuxp5e/kDxrfwOKjH8mOps1
cYPhCT3f/EFX920Qp9Mbgqt2vITKK98P6j/MKZW7M++pxTrpjw3Q4l8FD9dVj/xmLonIG/JwBUgB
0vL1VNQTjfvXpHxYmnwQ4IFZUeOvmzUovMubHr5p1FBny3B7cgrmIfYISgRhVeOqYwwAXd6XGG6r
MOlNPV/TkH3ndTEGWJLkOEK2M1f6eiQKlzEcQuJ0YhXw6Pxi5fNmHvDZCCgQ9nE/n1o209BGrcex
Um0g0j3oeuTvfndbuBnwNaFnR249rxh8Og3fDjmv4NtRqG7MSpNaB2QPuPOKNO+5NOgnLmNJ2X5t
3Ily8/iMSdyGGlNfhprf/+f8T/Wg2YzmNzxjku2ovEJopgr43K+F2wUO39LCSxjIZjnP1CDuv2oe
snOiqPKztYQuYIdkKh88j80dOq4t0ot1FvdCLHKWG4VbiNCSN5Ya9FONP0nRtemVL+eRWOjLDnfU
LhpVZSrmz8YTUkjM1ZnhSKAeWTtmZFWHL/a/adxzOU4O8e8MaOzvcsVRjLzAyIzvuUSuwB1hEhOH
2NEkK+uTVIRwzG6uMHleSbfbHWSM2q1ZIvnxNFEbKOEijyOI73wEmnQgEi3hwydyU+UEFIq4lXrB
UA8yTTNcKdUuKNpaIvpb2N2Cz/CU+GMQ9x2suZ1qlV93z95jGVZ/Ltx2sPG6gcWjaGW7n4vZyElj
+P4JW9imNYpJKUNagck0u8QmPqPeBcwFstCflie1A0lr5BF6kxKN5ZlbYNxkNymyJuFlJkSSvraW
xC2rfHXoL9glZ9WSU+3nv0tEw58g4wrn4S0gdVLfUbx3k2nreTe/tG+JGRiMvLpa7ixk/JL9m63v
i/BySNRHEMo8lg+n2QbKSua/bZ3PCt/RAUwtxMKXgj9IX1gsWSzWytUjom/FF87iZQCDVfbvjnR+
ifwkuoQqxO78lLGoIBFzi9QxoR8RACydNgfMH8AdYAl7OvfqWb1A44FfHUrGJbRaWhsN//6rFLC1
xUp7t7wBufyLob6F8JLLd0ZB7B2bRjIEz3mhKty/teo/7/sUCUp9hrAgTvuUaaubaexAmzh/5C0q
mbypWHt9alG2h1w5Jc5vVwTxI08d8cIDeoViOOlgHDnUVT+WdIzsHO0fCHu8Y1DXAQWUYTwl5L6S
u4hY+BiYIqF49Msfmwy/7caPiRwErQ8Zg36WbqFBlnizoLnLP3wFZY2QNBS34asIilGiJ50aKJ7w
P/oKRYNW2oe4AOLgfaZ29TVpibL+dcwxVP+Tgoa7qfhGIUzOXp2sBQsbxuJx027eUv1UdliEJjZn
PhDDwTGvRYONVDZ3a4nh+VeuD6vZniVJFjLu25zKB5RNPmS/6ZPC16qCRLryp5mTLhSqnXQFrbEz
SrrWKymDmqi6Y267swgY/0KvB24mGq/xpiHQ68jTRmrwDEUMDlPielB3fTC8cwmr7LULzB2o0ViC
WNYrpx7jTE+PQkeKld5Myo0bzsszwALETKC3OlxSfn4NGnxemV8xShAD61hFI4pEkaMrZ+W3ahDk
b8r5H43d3LnEZVZm0CDerM7Vy08wJ9pRruAXUkqnJvStEZgdkcsb9NLajdaiMC2zMLQ3AqnKbFz7
5KtrJ4IfImeE2QNYxW9ig1N+obS09DiAjHUMY4Aw8Ka2PFJ3fSJg5FLLz8U3EW2iJnZzJD8y389A
9lSSyyT9PF5rrw6BPOsQ0LquMWkNzsohFtfTAw4gnwI3pxgaEaTr323XSN5H/87FnFUxufcyTlwW
qwWZeM4pIAoaa4A1Lr5iZYsrsp30DWkOr2bgfXEvEGoElR8OaPWiHV0GQ5jxu6hykSLFCfajdLII
CQmHQaerWaG523V3Bb24qyOiWpZNa+jwysG3LeMdJUyv15GNVArv/ElGj7CQi/e1zfO7ZZaAmrXU
gEwv2sGV/Mra0CkaCyycOWhps9yopCbfnGBp8l9A4JXqT+bJGu+5cxx9KLiL7fp/qKk5wA8VO/al
u5NFME7+EdVn8c0vjhH4ISEn3pASGYOiOK2bFMSvXkIvMeifmA7v/NNqQAZSzGDCKb9hAVgk87p6
5HeThyCcpCeogF/QegmmnSFLWp+j2Rv4wym7lFGaUdfNBYVFtlkQaLwcYylu72vkN/+kUhQZy80j
LK6ccVODeVTqN0SZEkBbMVR4qAzubx8s31Va0gLh1qfa459D4dOsqqyMB0cU9c61evVxtFQFNDCT
VRRSpbWS0qpwJgLSgKq7D4yHdO2QbfYj6VL0KSSjAOJ2F6dKlWKGz2UnDkI+goJ887TPSmsEHQOX
h3JIiSV8lUYqgzW/IWK3kI5d3qeb85ml8drk6z68L8fQg/AGtdqJv+u8/H7o6iMB2pen7bh5O4fc
moYjTkjVCokdO/xxXsIHCsgiFwpaepEJ0plM27Z3j7rRSUShfKD97pKXt4UCjbNx5m/5AqpchN5Y
G/K1EHmpBf28eyp3SImO+2apacixBptGMLQ6f5gWDerNT5ox78jexjGVvXAlf3COmt7buMjGxPPc
Hbn7Z7Ps2AmmnkvNwb5SRdJ4JfAM9w7e/d82b/1/U98QDRtY/9piBTVeROe9QW3SMG/J39bm8kzk
zIjrWSG1Vg1HgSViF8wel9XYBu+hAmUiHLd9wEzhtpBDMxYTOb5GH4i/Vaw2cQC3uCJFMYfrwVi1
gQIxIuYJZYBbIAisAxXE1vM/+KsTnUhjjt8ED09MWVixDL/eFevXbPVbQ2o3wsSlnJg26PsXTJxE
o/O73rGf/pGlgsVwer3xl9g/VlYHedjd1c7j/EezyftKvWVQMt+GQvRwTOODf3rArtHuuaZUbm/s
yhtQYUhTEQvZGS0ut+CSf/mWjmy/0ZPr/kYTIAdDkY1fj5Xcb8cHBApv97kIKCX4GAd+xxckARQo
wzFyk7DAAgK3EpQC8tP253s9K02TmBouF91JyB2UzbqUMegCQrL7EPBjQlU+NXPF9Xmw7HMZ86LA
GUEHalV115+H/bmqqkuJVpQiLaEueV/r4f7qYn2vRDV6955akI/hCcW2WHPESie1hDJRhKvYcRCG
v+NCVur1cC5svZDoSe6FiZj1Xs0rxqr8wD0Jw+dhS+klVujyYLJkXMNiiki/mGo3XuIQzuvDTWeG
SJatF4c6NZ7KhJVfmqft/6/OAuqD6SG2W8yDJawtNKGJuO3dxjSqv3RO52xUgDSXDghhy2a6iZ6K
kuHZYrYF3VsRahv00o/BjWs2U69MDzlFeyXzQmLFORsg6FuxuR3zQEcAoGax88xdT5OeG8ezWRRk
jgxRsuM9i41qXkVBAiYu4hHQ03W2v2ve+2kz/Uzaux66sL5OTuZ1S7Y53l7EhLgHIt2NRuq3VE09
ZV/25/M1xYr5NCZ7PNsNMKHD7ajFRh1ZBElXVM3wPli+gm/npcRt6hCkCyrniqm87cNTP+hE9zzy
EWw0vAu+KmTwRhk/A4Mk9rVlV/s5gMUDQDCaivJ4jbP/fdybo0NNNxxl3Hcewm1zicgfuKPfzFiW
SRIxwupZ3WpzEVSUSUM7BV1PyupPZ4jlHzomz+FuZuacB1QOw6X4DPtkAXedNn7xAjjkSE77yYog
M0hpYwnxCWrr7eZZ9TsymVGCy2anxWwqapxA0LLe9o2McP8+w5ZZxC1nVfCZ4QiEgkgY+i6ypNj9
xqLLfEPu8Dz9E/QXNLwziBCHS9EyxROaScRs2jhz5UGUmAikpped7rAYV4a4eq1rtUfJzaUv7P6x
DUXtlBIy4ZkZPgf/ZK9jVdRF7zhs8GOdBNxLxbkUJxHfhT/Ayg11umpNcctdZ4rjWjqZKjS+GnAH
PR4l90vfmnSkHuhxFNmfEKbeEIUk2jcYxkVUv+dmAt2KI1CyQ7PV1nRrpXvq8wpTBIqowuePCPkl
vde4l7B2qfvNUCWKV6FboP/76wbZLyagnYzay++6ZfGFnHDqam+mhD1rm3QEROMPWj+CTMNZRyf2
jPz08dv5Ag4b4qfu3eNCSci0uUntAjlG/hRLK4TGa2yU6OwF2agaIZYKlwILLHRGylR8/hVUHHp5
qqtUb+4BakdPjN/ijUP4WetT6ZaytRKps8ZhBjwtyC/7YjRRCohV+1nOHbQ4aqwAZNRn5LmqXE0P
F0MyERVznQXu684v92ht8uGuImcmHtGMmL+EZh+AQXUIIzceWJR6tWfQZCkwaWOd0VlePhk3wknu
dBOmjzTXUIEni+qI0RAxVcCXNsbmPePu7ol68Vh80ghqhJL+HrqiTh3dNZ0UagH0DxmMHspeei//
y8g63ZGmakpnmrv/j99H6H37bKjpyXVif9MzapiS4I7Pq2aWPnyYdBGQcqfDH4KFhYzY5E5kOG1o
PeOFdmpziqPQcceuFD+pAYqx8CUyZ6wcARZ/sWiYJ4wBdjHPr2Rdk2ZGFipuFl8FYkiivTLCmENN
zwGrHbJ/wYroYgEuzsaQcmzvCa/P6KjKovjPdj9MkXt2GHY+detCIfPrGFvwroqlJbU/4H6fhuVG
LmaEf5HQ124+d+/JfCgopmy6Wi0Eb9H24YtOkH/HxRwYUcHbR8apOXsQj0xC7WlMQE/ycidtQhiL
bf5MeYQG/o4UXpnztv78YOrbkXp24ZpwQZgM9k2kvii3G684QMXoskZ0ca/4mBIg/egH2Q0cUsHp
A81P4F9qBw+K/tjKIfs2+1yImA0DsANBiMGJCB+Syn56i6NOti1ANi43vIQ6j35U5S3rF3nsUMu3
3uZ8wsBGpOa2tz6OmCSYEyNLZGPUapfa96MD9KxpL+t3ko3cHT29fySFOzveVLQ2COWbbJqFvGfl
LziJwvpGbnTxoO9jBc4BtImI964mDa2gZ4TwDA5qoJ+gDrAu5cYrPywTozyBUvSoqr63vDTGC3Qh
0pg+6HZAVTw39gfMvLbK9hiEv5kD5CEjM5H95Y4EtW0tRIqyYXIBxc42JC3OOFro4hEPAJRChE0i
eR5qQsrSJVYrFtdwkfgny471p4UYo5nbgH8Kg+fDPjzZRwl57DNsLvAaUea4B1oHbLNawpIGSfax
fT6TKvJygZafP1SWyrl5DCCiifF4C75uGtR1F48HdelWurbUkEIrXreZUA2og3n4pHu8e3rU/Gzk
xyUZqcExwpupPfFRBhYbiZ9sDlzFckG9HIdRwKtGjlQrVsPpvV8gsAEQOsJM+SKn6sB4Yhn+1qAG
0OcT3rWY+T8m/OrwVMvS3ihcN4XXJwH2jGw8uuBkChzqUkBhQGXLZx+wLW6nM4JU9NKzu9BgsYes
EbPy1Uph1BOkWLGIdZNwqOO2Uqx/1ODw0eA4f28Je0ndmQEBKc9p6Y1tIgdXUZl9qZi+jxv8UuaW
BHZT2wtbkhXdXNbdu3uCqszqsSjyax+8LO517irQ0eKYW42o/oT/LzzQ94rSXlHvv9UiB2geDEeE
QcE1o7saLcK316BkZvUovIkJL+ssjpjupvkaEIvcVBpQYguBcMSaSPPEn6bquAG3R/3xS0OAhwTq
AMBaZOzoLMP73Z8xGlQ3AKWbEXupsD/2OEprSAkEhiJtc2d1v6E+2QellwFm/5bsAKIVYFNOnLV1
NEExGqIxbT20uFVI8ebLEYvcUFVd+0zhTJeISSD0LVs5iT+7xKAWb5beoGMoGPZLNx/i6CVowXGV
JTONk9XKj4iENQpcQdUSJGLG5VxTM5Zh/8MisKbX6pzXB7gQ/7HwxhvD8AAmFx7DbbAfVkryAvKq
/FDcf5u4VKz//hznP4el/KsrGBq24jMIeCU534qgukb1JnUGTB1HYorgMRA9+TPNqfF9KTAXkInI
zb6MjfBvsiwsLIzzKbyWfNTImYEjLGbB6gVRxAGRg9+VxwSf9jYxhG6iLMxqTOqWBVxsn6ZbZgSU
RKVrH3kyV7AWTGpmWpkjDnVYQXuQMZOudO2NXRPFCUE7MA39liLkPIz5M7D53Y83+tE79SVG8ltP
i+Emx5JgbaLoysafGtERDM2KtqGY7U4lt3t3odTtz6yJ8Ol/a/qcqb1aBwrXer+BTL90iXvxOkDr
syGm6KTW+9vUN9gGx0NVZGO9Ci3XuqJwdoM5zy71qZ21OKQ1qx9DNFFRqSaSkdSuhqzc3euUDGaE
3DSM7r4WBAzR+7QXOJ6hcEtQP42RL+P/uAYjjIw3qMQSSUNMpZYcdbWubV+/Diea9iCLEGhPBKgI
9Ftv8By/HKqy/wyXdper1sbPwCB/i+uj67XbWFYFb767VuWn82I4RzVw9UBxGxvv1lbUpKPCcrgP
XN3RObfWc5knVS6bX49DSQob8qn5yY8QCSzmyPr9J7YsAQdyYrR5d4AW5lC8uqv8bb/+53yeNS/l
Z5/PRrdg3mZlWp3nCfI/6M78x4Whm5bvakgd3gxiigm9mzn0GlMowXNLYx0fkvZEhPq2iWyn5gTM
/ul4b4VlR28DagkeIrJnCGyMxlGtLc1Rlj9p0SdTRsilJDmJdicgL9tw619kaiA7zbJrIxKhvGQc
YNQ02ErCefbn5yMdlmsr7k1BIiE3V5MjUG4nb5TRADc73hD8Q0BFLDCJbJchTslj2UuMJEiDO29U
YJ+ZqFbRILQBJIK5xXox1U1FduAEh0f3cpDRjlBvE6EZqNi6/97EKFyFNumobO6IxjYyH0k+DK5e
MiOp58jFMDd3uLPFEQrg02yTkmZh7BE+smm/kVk849VCS7lb+qRsmtBqMyTtI8ezEsAu/STZY75a
NiaE4+Gph50OR4q07nBBPGNX5ZZwZY3ns7pRAnroQXJcBu1WTuz5K7JEngpE7wYYxfhsLVcICoYI
zs/wFYT16U19QvC+VmTX/gfMysCQIvLxIs4GJLUGxKQXIyp1Gw2WclB1bnsEeQEFkGi8OouhIsq+
9pIe7nGtbHQoi0ZGAtVrx/FPXewj0i51eEkQQWFkSML36cU1ickdDxJlRizEbWspxG7vrdixRVLZ
U+XQS9mQV9wRtT+AExhxS3M4p4TyCtnrX5hezn9ffqoXjM0u+SsW7MJg9XhsuO4/5xprWN0S3PsR
zE+R18rDgpdEi7Dpn1byw2wFmCcPl/Zn/mHl+yes6XhUJuyd0Wb4ECeR1Rt3UOYOT55VouNqob64
FBt/qSWb2arm0CfnlAuxuLh79o07x5pY3z1sJqr7jB6s3H7QEQClv5ZNcWqni4oXUQuymcDtKwRF
5HntR+drSEZFQG5X77FefCTBhZJWJtVPDIiXfZcMieVUJXTev4aa+sB3PLLK66pbb9zRu/yYiTji
Gzow7X06C27YDvICkgdg4DqF3awqQ5T2gM2vAu8DkafwYWiinBuo+PmdkntNOzDJXSjGN8k/bnw1
abYvr5eTZPQuCOyY6qlnrhSywIJCFDUVIDgXZRy5jpvNTmvi2vb+wjt6Yu8lS7eIzshxFPD8CiOE
r2JVxcsuCkFgbJoweFxZLAsOsWxiw0rAXQNpnpU6gY+RliBI/yZETCStxK5RSeUg+No3vdkc02pI
JYzlQ+a7YYw8rVDU2eWQ2xtPyTxZLny3N/3XEQa9ZoGnkP93TPBjgkGe0P9KFopXWA5n1+X0CqWZ
892gt2ZVKRywh4mnaG1nMgHaYECLOh8+ZNmM1U7ua/Ta4yB13e0WqYytsSgZIDoDz4MhG6ZWdy0a
XAvcEkzw1c4hLOFap83pvl2ID5t8PYa+Sq4SXucUzrqlA6O5C8gqRXebETSnrIVVX20PscMl9W+W
stzO/HEb3lM1HPx1xr2HZPm/0Mn0N+b9LxK1w8ThpEBm7JVaDqXCG8M7HqjvACybtqa6CiCGdGRE
VFacNlj/GPeutDkXLNM3l0/4r81KEbYWWQCZrR1ehJcTFWjMuA3x+TcLUODN+KwN0KRu0y3Smmk1
cENcUlJc/E5PVsBj+LSbQlO37Wo7/gkDcBJIKDdagwltqbJX8dv3DttA/Q47PY0KQLhHAhbcCE9L
KKoSfG3GCC8tvSk91UaaCRF16JNGgQsiUj4L8JFoZ6ttE8js1Cs22C8ftly5bjHVNIepkOXqA2G4
zORyN7/c55HHZRdDsMNzORGxAPA0PrZoN/XiAckqWWiUxaVJNQ7onRcCfrYAmILTkv0XjyH+qnUx
pPwSwjveXivxHSb/TLVZbX4O2rylpnS8rt1sV3C2x7VIdbudCS4rp47q2NYlQAiSOhiGIB5g6Qup
pF4bKnxL5dZUDcldxCpZfnB+nZcCaT2Br3Awkx+1MU2vmpzSz005L1EaZbiyIX/yWtAU69LQ2Eqv
MVr2zeJVWzRz3NyLuuuV56ypZ6GrlA9yOsnjg/gC+BiVOWFmwu9JeCAcKiYGD1hj7mnb+VNIWQ01
MIagB4Tpewl3Ppdx96PSBFOeXpm9lXYXKLFSsVA1Rugl24lk/r4dgrfF2boknTu0G9HXlDnkUFBP
is6x+k5pEPkAmyxgqbuQ3dA20Cv8qdMXuvUMFSKgqvQKQz5GWxDmQGbKuOPmN9RT94THeXtPj8/b
OE6EmtXsiVB69og1unrDMxJwq1mn9gC49w45M5MM6pnAxvDMQh6oj4uYmM2QxIfw2RuPVoIZDGLL
3djInLg6mx9oyj4vG5K8Wmm99Zp4VpJkSoQWDiyZMo5DtOf0vDlh13So6Cn0nJQyoYbcBq/qjvre
5mJjv/zmvq/yWnnF5u0IZV4aKs6FR15S+pw6m5y94OQue2Nk7zveAyEyT0EUFtvjUzl6MtggsBO1
CDP34D1MUlz1E18M+GO7P95Gvazsma5NeFayy66WqxkVTrIpA0kelW2LMqGgaCUHM3kqImKsXDDS
cWcQtoZ9t8ltxT+uRvZrwFQ0y/TpH7F3xb0zbFXWst0Bv2lOsXCCP4Rup0nCP+GKhz7mkf/QUs71
vAcqiDDF3D7seNQXIC4NLgB7biVjppnBh/ANIecycF2sfBOwPSUM7wV/HsCyjYhZQO3RknUec7cF
/RI7GaeWa1BPxQE1BKmsky4+BvKlxDt5SPXamjB+hPeaUQWwPBGYE5UHZyY/ePV33No0nsaIP2t2
wnWdtPGpYA4re6Tf/fTGTJZu9pYkQw9fYT6YwS6bp0oZ3M3fOw3YzOKbk4WfP0GktYwO8ZD+2QlU
Cz8M7swiQVNhFQC8O8CJqysL0VP+VlAfSYtBZpsa5ruQvoZDYgK2WESdFZDOFdL0wXMcidzZYw6x
VLrPZMo7U6K0Erym3L7kyEneZivzADNUAvTN4YrGAeJRd0qbFoPikbeC3wYauWaMaO+murDFkINd
XrK9rzdYJ44yfYR/h7LfZDdJu5W7pgJekzS36EDk6wjGZSrhNWXxqoMJyRmO4WN/ObBSb8uK6Oyz
3YOpgbVLX8XyKs4TEFFVzMNzjraJlz0v1TsCMdbMafVb5YeQEHqCHkn1zCiCn6EEWMyAw0J3+KEQ
ZqJdqc5deey4w1e06Ovsq1wWNPbwkIfhuzcUZx4zKQtXKuBH1fL6VBgjGXJ2kiqJ+YdteYpHoikX
CpXyXjRktwyurdH3ArFrQJUZwWVHK+QDAnj9Oq+WBo2dMRzMO4kNtIYDXP+RkFyyywlIwYWl4XQr
jMr/L3t9enRM+fY6/302Yb72Tse050a/HWuPSnH6AlVEig6rS2RPnqcok8ymlqjmf4+AgZ8RKOiD
nnPkR4PWoQJ36kHOh2VrcX2AbDdVcHc9g8ye2Kc47/yX0rH78HYEovsg8+GgtE72N450n5gDF2ah
9GwSgpp2PAHTFNcPxNyRz7klZr/jNTZ3CrAEYj09oZs89eSx6+zZzndD3sx6i4PTMfqT1Oc3mB2X
EuNN0Cr5ZBhjmfWGLCcCTeuwLZOQQ9tSsdadKHV5ciEN9ACVY3xEaIrtExqzTsySOERsdiTZS+mU
k0hmDp+FjeKBOjAjSfn8i9n7noHavf/mHrFd1WJPF9jYvew6wP+GWsLZLX6nOKyLLY+2cY/5Ie7c
WE2AEOLfBBzMAfo9n0WJj0syUbnuSeM8HPkStpskJzJsY4Juo4VAuHjr0qs5cSnVr6XoCF7cXu0p
zBIQvUmVVFkVRZiWdzQVH7RKlRQvEe15HzveqWh+BJFqoeybowZbgSLOret2mSc/6V0ul5g4QeIr
2q8XJeoChio619vJtJyRD/s0aiRB2KjH2T9Y30U2FytLmlVU7/tyZvxk/e4cjqdu0P01+K6oSpzd
ZPeLR8Ndv2ykhw1CTaEMeoFsy8oXVvJELF5mYAr/rkVLw7z1kN1ilhnkdWKG5uFh7Ni4hDfo50bG
x9vjp4MB/YEBer/e9LVnD2q5Ba/gLPUmXVoUvI9GVhOfWb2H+L0uJCAEFyvwR1bQRAxj4/Lus3q8
h5D2cbdnhEIsmYGytO5xe4gqGNRvVHF5EXdSsYnLS01Ahqm7vVvwFPtVZDx6jisfN8iJmJ4tNSeo
OH3xzwm0Ok+liNJnXVlmXYfkOeZKybWi1cLAuMbnZn/W0VXXbHX/mkg7bSUxAfSSJy8t9KMlLcpD
TMeGpG7ustUjkzfmlJ2CCJVUmZJU12ezfHpv3qQ86e0D41XOI9T8zPZqqRt1b+t6oUbIH9ngvuHz
azPXeSACj9EojrMWlI0sZnPqUp/ufFKBitV1LXWs515B7a3YT93yUSZ5XBT+rBcNtM5qBIJmI44a
93GEIePmE1nc4VS5+wT289Wv7I8EEqNrGC7Eje9DMxlgJsK/mYwo0sunBhaFhwIj5I932lwjxIa3
eoagTGDoseGFlreqAsFgFA99yYTj52Ang5S7CEVHeBbkhyMv/Bf9aJKpXuF/wpXppSYW5izDLKnP
A1RUluI4K0KzSShYWveVRV1VkeZfXGHwn7Xj2XYGZxWvl/+9CByrpuwGiTwcuWsa41ICDWZERHWJ
ng46XdEJsbJysq/saOXOSSh0LZ/+F31dXuCwLQisc6RmbOlsfnW9BcDYVZN8GH7PHvrZjC2nUqls
kFJE8JviIKsC9JdDSnnyxxkJWA5F5Ln6LpnXoBUgmoA/+Cb2WzLGfrTaew7Nyp5gbIOjW62Ux9NE
Y21w0qUCpxFGANfIgzoDhykzNTWUAXdZd5CF/HugUWluV23hFTNYCEaA/hcHky3Hxad4wsZXIEzM
yKZFhvuwEvRqPvga4Eg/BOigc5vVqSU9EG/X+bbRpYkJUWnWrk21iaVJi+ucHTEtK79KRN8pQInV
XrFBuaneAkyu7xwUPFgg8nJNy3PMq8fcaSKqrgHbL3sBAj/fEqjK9knpb1wIi5eeQIpG6bqkXdPl
361kTbAHQQZ076ibu9ZM/yZTyPPFrocKAx/Ind1T1aNlK8HPm2/so1rrdySc0dhx4WRkzMDMwWv5
m15AP5m9ePFUnCgNwKLAmQSY1weAzK5YaM8ywaBzBQIiRFkG9YldIayOp6rUxKKly5hgn1hCZ7nJ
bnToAMr9Zibl0TqFLT2Tm1H3PTV8q+sarg2S21PVd/WWu89qvtc3ichnoQnuvwdH9+VhTcFnvRnq
/MeC5Q3Y/e2vejxgdpY6+NXtQ+VbzKawro9fWVBgCUEtZAEKZaA7CT6pvVUIogPwUL6fIUqlpexY
apvTN0ngUJHvoXvJhD0UIOEfyHBqJ5sSiWuTr8OoovqbthkCVN3jRsKHRB57ZZE/DzIUkF/cVTi4
JULwAzyrJkdGF149bgnEcCsDFh+uaDAfSxQ0Oip7hidKejgbukIeOYUMJ30A3XbFQUc6qQ37Jvtq
sfLqp6VwKENw1mbTANYTOw8tc+8UpJ9dbpoNPSTVyryjxHY+F7oUttyxp7VJdADSRZd+ZKZom9CG
Vwbc3qr01gPjFkalQvevu+i/tJkP5YCM+go9uPZkF5t0lhtalGK+53fcwrbXllf2lDVINwr/R6Di
rtWBJqeZIpx3crVT0gGQle0EjpsCb2SUxoeJ8UpgXDn8HDGZmMulX/pSkcHeQX3R5154S/qvF2QZ
WxuQgPpObrvtG15B/1Ui5g+NQA9QG3pbWxnxTthxPw7pU0lH4dFV4A6kozLaWzJAE3wrZenNnYws
q/yNjUbMwlTf93soBE5O3Yu4J1aBKUJxk8nYWMCVjcIMLXLbI2uysHHgA+GwaooqFUz1LJ07bdvZ
zCTydK7T8zhkpFbLixt9uAQLZI+09jpRvDY6IwlnUwieGBVAZCNlo3kUrosE1zYlNtLkycWjrFT5
jU/Euev4oq8cS+zIygrj02AmE7TRcS1sJRywaTznYuEZla8eBd5jTtnj3JN8rHH1nX2bGB2FbuYw
JnxUX+ocTY7OE2I3TcQyABKnS/ZCIY8Oo+xmNaiPrGkyAC7YST2HKPpA8uFt1l6Ke60/sIFjnOOC
FXMcXN0UH1z1e3j7BCP+1GR8gGGzWGSIm9uC4HuuLAQLJeHcG+ygWt7bxGCg2JIfExUcA3lc25xs
0URlHFxFvtIKyQcGVt+g8k9QxIx+M82UJCNBEs5pGKj9BJqQTTwnD8B216pH7Ze463qlgnMm0Plc
sewQAFs2gjH4bWH4euMmZYG0WwWJl9PI66QHvoUK1ANL+f6XYWB34rg7sWQUFkSyNNKcRyi9gxDE
zyZVwZ75wifQLdhp2ZlQNt1A71kfR5ojdUWD2nVYkzs9cNJNNagQw5SgxbCSNMg9gvWg9mkuyhX0
jugNMvUE3Hfd8C9lFBmoexTW3snoDML2k2rXi+b5p6yds/oHpSZPHvYspVmWe7AUe53z+o1Epydg
ZaFDUobi3vysb0n77iiP4joMSeU7UnUp+fdCCqv7y5otZqcwfwFWPkx+VuZzi+yQEyOwCuedJx+y
T9wUP0bdKTpqEBkiBMrjbADo5Hbu026ngLEGdNjG/4vX5XUMmXEY0eQ/CqG6XTLYev95ixx8IMud
+LLIyXmokH77hSdrh7uvCPsd4e4MuGRN0xjCjIPypCsQG5rQLbYWjqQjGnRdnzUrrErRpwgTRpFH
xc1Srqm0yjancJ0EtVBzTCUc1nAQY211xLdiNbMPLSbO0YkNeUP76NT2HeqUffP85mQffjkK1Uv+
Uqhys7fC6+HQh8BJQHNmPJqLyyqscxXc8v0Lio+/hF1UN2CtKJIxh9m8L2isozMnYD/qAIchp16g
UUFZ1b2FpW5uTt//nOqQ5Aip1CpOeZWeDskrGGT/kvs7IX/jRCu3dKGkiHUwuIoRzyB9KVpci43n
y0sA/MD3zWEQEbf3TJUOT0uakECRgHf/zMgG+YxEZ919lccdjAEl/SDwTaUO0SPOeHysSWqN5tc1
oRc1FbKehuJSF2/9PwInEcyCb+DU4Kmhe6bXmH9Bmv94xfEJ9VRowApckPBtYo+Afm6g22QdxNgj
5TCukV8Ebn5m/pBX/s0pbHOavHFSeP2Xzhs0Bane5uDb3VbzCnuaekvGwtk3wp6/FG7emmGPOMWI
UTh0t5iNuGUmRxW9QW4xwjSVgAOF37a9ipjIjduisH/LNJsYF3IpqpRGE0s+6c93W4K9Rb11wyZI
mqSAHTQekJDarTEjdSD58vhGM4BoVA2Kk6YvOPOd8M5JZ+KxhoDbN2pR9W4n3FoHk04EWWyyolg6
ibToTyyGZmXNLsoGVFIwvjpxxt5nrynATMGo4n75INiZJFo6Pk0V+Fax5CcksDO+iqOmoD65OpH8
6oHiQVz3HXwDAQv0O+ivUZc0R78fnQlDGsWCoTwsmOpSo2bTw5+1KvfTLkZbwWd3qTKTTnAYtQ/C
V/Hp/obLTyJLpxfO6OgW+Yg7wgjQpJAs502V0PWwucsG+m3l1tPzgXT8LhQRi8kFeGaWrejZa9aU
0OggSjgXWsJ4kNqK6w3smHDj4FdCjXpPWW5ltowFlSrhK/FRgBalswDhxC7KKKLHkwGJ42ZhM6Cc
tjybPVDxs5osSGwYq9o7yqQGmPZb2rU+Mu+sApQvRRFQZVB+3kjPyyEByzFIN8lm2sVX66+Lj1ry
So3VfwqdKteiNWXHADczKScM8Loc5mS1XE10Dl/Fg/gIbzQG2t/ihaDjTZ66Qv8yKEI5o0BdajBK
TuliWXlqIeqZwHZoSqFVDdgzj4OILB5oGgfLzfPU0d2PweFwDuNiyvzG1q/ZQsxhLbAi7sgO9BvA
acmcY8Z+u3ueZTxr0YFYc8AdlbiAq3gGxhQSnMZWp/SM+pqnpqxNyAQA1byV6UPxHtl48+71J3WL
CNNJ94jB843OhXYfoM7MPE5tgREMcAsb4Zsx8Q8AEfw9jH6PPLpazajIehjWYNpCwmTIw8WwrObV
nl/+oLL0oUofdgdSkT781NtvGSwJNfpfnDWCx+TK/F+SdJ/ga4o74D3nm3B0qSIwdf5nla/n2+LL
pVCIpsZc3HdZRN21uRUKym2a1onyZebOZbCBi3RTGC7n98wsf7qVwGL64L+q04Qu1InGZJ0lEXNO
rvFHDlK10YxzbSvsZevtEgFjimNnd4+XD+9JM1YatwTBzNIJT/17tdDhqNJaE3JIO/pIRfMLvxDE
mMXeNQoSSXwOHQ0abLUZhJel2oHCkme7hvD06H5loWQqWWu3ahX+S4T2fUT7BR0LitDjmTQWR/7k
u++tmeASERPPy+MtlDeb7SXDynnmStvGHASl5ZxCE3lDOdwsakiksV4CyITVtm4/fjn9kjd9ePSx
EyTayTEyY1+4Iifcoqyy3h0pIl8ev3hKRJh3akFDsUm65rtS7eiJ0WuOPAA4QzkWcXP6qZ8LHcBY
3E4zZjlyUqmZhsmUN3XOnyr3oF6Vn000TI6Re+VDiK0dXMJqdEXafydQ/0NDdO0b2wuVcLuwFDbL
6N9KTIqZyVuGPxh686h8HYOfTdCQAJsAuDiry3e/srD2nctpvkSdBj+9pnZ8ntRKImjJL7a4R1zf
RSUzqhOlpYDG4iLV+h57B2EjHrTxohHr1NofldSJ2WFbSo9Haww83TvO0YWBVXW/1awoFaJnpr2m
pX55IGaqip2y8wdu/5gXjnu9sQiDXQfMxmkfDPUdi1dhRjl/oiw74asvFoIg+jyFtPWKllKtQcGt
11Tszbxyout5XSa7eh0rgoaSQbRegR99pdJ9Df/B7JIfb3hkOvqrpZ2/4Ts5RbsjLSSOQaTli0yL
HZBnJhRpAJqispLJjZBbcQc4z/vjzz8rtjOo4Mgg0DPZRWb9uRGh8CQ7TxgAqs6OPw5J5PZYpJuO
83OsGzfkn6mvN+gqhx6nxWvz/W0niQcR6QzPMd/agIoN5tqMYmWzJTJgRsD/0ECso9KpB/zqndEv
J3sFBkUNZlq7ZJmYvFfbtH3Bisxi913AcSV2E7iheFPDFp6LAn+2Mp9VcKyLLMQys6PqT5o0fNn2
z3SKErxbHahw8JjKAlx+idCJep0UhDRB5GjT/DeRIayKr53mu6S3UQleqFixl8vH7vk166qe9fdK
yQxfCvehX6ANTdcjBwfEZDg++ojddM8gGWFoHf7NLuTPq88vb5tCiigGp9VqM6dqSpnRvOgMXzg0
JpyAWn3DNI3QYRtw9DqIYYv0+iV5qbyLWkfN+x/Ut1dJWQHCqAc56YiAXnZF7PHJagmfoWCTo36O
niGeSaEt8EGZVa5Qfkr8mybKrb9MLpi/iC5trylVobAI4ar70NGhefl7gEFlcTAHfG8mcUJPUlVw
gUoERev9nXYIcU+eVxVzeOrWRVWd6AUYhWCDMHfL5EyNRG/uDKCGGQh5ngAdq8r8/M5q5f0TQ/r/
LCgbYRAlXTKIkUXjyll8u+YbjwcUw2mBNgPo8X+GrXrV+3O6VhuXMab4V6zN0Q/FX4mE/luLwykn
e7clC9j0hH/sH4IzLDvVKgrhy8Aj7csSnvJucYBjx9r2Y7lMLPcRuOIvsvv6SAQrYzqT3sEDdRUE
+dZaA8CGj0w+BQ/mQbcEQ/lQRTgDNGkowipphAWfdCe8b8KWSnVjnZXKkMyUbm1uWf6YMrrIpzV3
sclvjqoO2mybM72CQhc902JIPsZFbcDYpHXl4ifSkkQLt84mejf6VG7wLcgxOYYZmu6bWV0zaRT3
87nC76A+Lh62iMojEFXtuPES2/JyQ7t5okEfWrIan0l2IAhy4FAE0HaCDECIaY+bG1o73s1nIaQ+
YcDdVuoKb9P9LUTPm1IbzK+GdaNmO6DyPyCGL4g3YLRAyCydHFxx59dJB75fgn6lvhdEjDbTMFm3
71P82l92skEdoFPlQwntx5+VnI7/4anWLyJApb4oAujiE7uK+b24AhvzekcbSg6Sbx3yOiV6U2nu
/6z9bgt9fCYgWhXmnz4Q6seRRD3/KBWWXVc76u96mmqr3o5MiC3WYiXRQcx+WfnHP1lDDddIVN/i
u/Z0rddO6sgpCHNlbNCslYKgwrVuOu5djaQn+TAfwKpbMFlw7v5Xriwznt1DAU8OeKEQLsNP8h5V
RJdT4R+ceoKE0BwViSWSQq9G08422S9piyyB/lNU0NTcgxJVmopiEOs0R6G93kaB6itOQBWm4FJY
+RtFgKgKk+RLu2L9XScgRLM02hqh+glB9J1wsSliQ8xjeEcnA67k5j+sbQs48ebvtR6mUOwqXJo0
EkYHPQDEEnfftqOi7c8QTcCZWWMvRY8lUaFk8P+cFjw4SWALVPK3slDwKUtEmAKpiYLf3hOdblcN
xxj1YAJ1K3KrfnNZynwcT7SN3Vji4cL5MWtoJjx5dBJtCXvR/9wP4EXHyUcAucmUaHSctROKjU0+
Cq1xGxwSoj/qPlow0yP9bUEDuITSSz84JHHCwKW9MIsjqH/UvvdBrUoURJYoDRRDD6caPtcS0Y9g
QWFJACQ9W07iM1HVEEItiqz6pCgb8nOpn88K/g3ljeo+xZhuFb8gEZUmx08Oi9dBs6YTDWNn5Avf
/U3QuqBHVwdBoWAyCX00g3pb8+AtBKptkFiC5YW4nhPhNGLBmBl1hSjL2bGwktes0RaAJBDeDwEU
FtmPw37l/42EQv2kOE9vaayjvbxHzx/joYhOx87I4XO0UuCZE5Ur8SAe1gVX/a7RVUlqDA/8qro1
mma6OyANXGcsIjTkq89VckzBhHmUuk0RJwW1yFFu/E8x27UrbiWajsG3vGQXNN/CqP3qO3CKXQqy
qWqDUPsZDQYf9UcLgY9BbiN0Ao0PRkj2GYxEKh0kdBQYPMmN+EUwUG2DkDknwKXKUMAj5cFPZSum
cEH0kwI+9CiEBAteL77jNEfC3EAG41LzRMO6bXwMCaGMqdQ7l7vOuSZqGC4iNErrzOSVUrO0PVtl
wyc/cIK6DglvVLix8HE+xnjqEqdyv08j3Wg5WiDAK81dkw7fAU6e2iW5ezBAtnKy04WQi+B+dmJb
7RJNp0AG2CQlufi302snEXdB5GG0Z9cO7YBlVLzJikyyPwd7Fjuk7LqUqGTGqBeXVwtGupDchrfY
CE2KLkBlZVyzdnv0qwEDmQno/28XPuHsalKGMHdmQu8LMwkJ517SIEXW+eajfssdouODENmzoBR7
pkdFLbBp+KSPmL/SyuBXc2twoaEVx3ZR6JixEkCuPTRL+xF8WDyrSgLt8Lz1oTRLCGn966stfXqD
9XGj0NvQhsPTy45yzPeGWdCgLE1jXh/7hpPPtfqQj61e1Rmp4sa3Nc7DkA0FdmWOS62k0wTYvR1v
LY8Fx/zUS2HQD7LwYbUQQDhetIMe4vvXp7MMHoP82oVJIXmwVrR2nJ1Y+VHeUzK+2O/Bwia32Ma4
e1jhRxdSZ4du/CDebIu2v9vvGXT/UnV9BG7rTeWPGXMFbRwQTUafGj0NrN0iF9iGYx8B/OlFn/7U
wmOu/Df68IEnJJW3Iaq8DRyu7mCeVRT7x2IYykLCQ7FKATpZU58ubWSlaIW0YvMQETa+jUtB2K0F
7+m8N3dRq4C4bZRpyz1odu/tEO01j+lVyxQwPb9jdfX6KduceBSDa6HHIO61ZiqhNOVdPcJR33l1
fIwQ4z3Wk5MUDsUk+FiFilm6rJJ2K1fQdRlYrJ3U+OjqAZ2X8SibF+8OCeaaNC2ttKLyi7+5taeB
ICfWaZgF4OYNnql/0ht0C0xk7aHSUXuPiWI6eB5DOAV32A9429eI57m0IYiDNXs5pY9OkTHTNDns
vkaE2JxummY9TClHNc/W1WzLUK7PYQ7fZZ4d+QCy1yy+VyKngg03z2FasZ/pV7zhCmVN998iuTBq
jt+Q1NNX0I+TZ0Beyq2CsIqIPb5Nra9VR4OL4ygYFi/6lxb9CBmGpPWnVCGpPvSAwja4aKCaA1nW
zARlkHgXPvHdKumQwmTn5Y+pFfYYCzP7f91Z1dxrw7YFwXhEy7jgJmAC+GMNi1rfsCkxlQqoxdPy
/lPp1TPAEHTGXIHZTsOyld03wALjObMzfvONpwBJigWq8h/XJHRyBpOrTRtBbkQisqiInd7DFzVK
se6+jvZg6WFxdwMDVCViGEFO6NjOOy3py8xn/vpYwc3yg5natd50FHWHmLFWeYbeRdNH5sOpsXjV
SBvT7nLe3gwRSVib9Ve4vCOOfKNDvRUxWi6uW5u5c2J7vyFW+u7uwH8JU+d9HlLJ7KoRnbZOtyg7
Gq2lo4MJsnThUiiMoDsfukTsU7Tmps62N+rjJkm3h48yYz/Nt6fz+gIezIw75zPhDZU0iOYXAlst
dIczSJnm+wVFQF6Yvsd9RoKL2Vt0hzN1JPFk/9dpgN4sOO28uLSbwefp521NSSLo3qHYytK+jXM0
TR0UYc1/EFZ/Dng+zqftOHHerAIj02YPiZBmx5t29ozmXj4zAwXURtFn/gMlrA6QdqWdBn12agA3
+HvElDhpVZlUyJ+Dsh+NPKIP7olqj3lFsFbHpSA9SyJsHlGHc8Radcgj1OWET9S+LiNEPnoIJaEZ
bFf7cdOjHZHGwBkR4MKduOrU8sHEL/p6PY0Dj5t8mttsCNUytM8i0GSWkgjRIJfJ7cLuAvPmwsFb
pzmNeb4hg0dz93Bxi9I0vWoBxpD8JayuyVJfWJqsOJKX+m6VEDSa7yP+UQUCkQCh6Yds55dOL7tR
tYcoiCJnzvKVZVv9nRcp6lnkUk+dfdgPo0CcNeH7SNbrROAs86XpsprZ7hgOiEZpAvSWc2bqdcDX
qdfVOQRZkYUyVSbsUtuzrV/Pt23vVUW1sGaHr4JLcv3Cpn0Y5iA90bD6blfMnOSsBTDyXpb9eujW
oPyXbg7yP1qvvzj6OyyD334JQedFe7xbcjur+g6w/3DN8hzi1ui5azvMCF3HQk02tT4Msn/9nQXX
fI7iDOAgDrUxiMBq+Fl2+ZxoDid1Jx52qakWUFS6bNEKtfjl0begIcjdMZmzlyF60LRLEXJsd9Yz
3UDNd8SqJG+hAsinCBCROyRWUK3LJ0rYmNlg64qPLv5Ua43l1NqxN89cztVNA23Xfsmep27eByUq
wzUHlu24/G16oexjYeDB5BiYSzAxynLCXEOCHTJIjOALuYg0cMQHc/V7ck32JAeT6l9rHE8pP+Bo
Dwxv3lQMlICbhvNzr9uPO2Nsl3cD0ON7VyrjBKMOARPN3G5f53BfKpBEmr7j6rP9fdU4/ZIEVSRp
zFLmxUTfIiuipN3HDVmirJvLjvuQyBF3z1q9xgYgrIYLWjSm8groIK4IXiYa0Kxe7y769K5HtPxD
MTZgqN5L5usi7sUqu8GfUTfDw9UBJ0kZ4+VBgoDDLIOmWwFywnyIOa+OawyW6FxbLbUv9tAfD6oN
nY9RTrmwjAfBcGdLjl8Z0Xh4Y/Nwm7/KmpYbFL3oPOX0oSBFLEz4HrrnRhAR0OdylcdXHr91fHfa
pBfeqL/l4ngd9YL8GRbmlxWzfYRkzEmx5sSI7tdW+kOTLu9G+CbG6h6ptxlmp/t6kWwaGLCdnGeb
6gxWZGUMw8bXzMD3I8xX74283sDOtyCbLLbu6oXiawPJF8MHJqNQ1KSrAUBMAXomzPva1+Z72rEl
xpE8mGDxfL31mb3ighP5DRepTd6qVLw/Fe61zie02K+eQ2vNOJW7JOEhyNrw/f4cTPRovNLDhSxm
GMBnPp5+Efm678S5GkUj7xD0mQ5Sw90ZkRtFV0F0uP9lAEZMpnwAqZQs6fiqqK2q8ml2LPkE66Mv
DojsunO0wCl7QdfOFIzGCqd5NrXIRw8PoUHzz6q2kPjl310SBHeZYq83zDAV1dQJyE0k2er8j+x/
9SjHQreaN3qYwv7M2slPE5+aACst/vOOf1TfiTfZCG2FF2g1I5LZoJrJLmp0VP7qj00uwJb6VvuB
KWRWAwdTzJPKgP7tcetcdRlMHmLYrvZepEl+qMnjOSkok1vyIIC1lESrwYi+7mS7HGoexOsFacyi
/D+1vuX5EPGDsx8jB2tOjE2c1l6AYu/lIIOCN3+xz4ZUTjTJc1d1PzITWnWyl5eLw8/9UVlANjKi
5s0QxM0iwbxZpDduC7m53FtvExrUk4wzoLoYPBPpVsD5uS7fUBTeTECYkiKueNjqg2ozMkYI7622
qk9TOF19SB+TMwwqss0nGY4XbF3Zn9We61jDxCPXxzYQjppc2H6gLEyXFzqQ9k6s3q6jIk67xxY0
rn9y70Pxx0Y1bag8NpZIQn4zc4SGP2dLI+SKbbIMjOm5gvuuuVNJ6XHov3XDWS2cM/Yg7BLILKd9
dwCLy+eqECMkjoIpUdLM+gRfz3ADzcfesRha7Dk3CElGgUZWuY1eqyYo4gnqoBSJEtC7ELd52UCv
asiehRnfcBudunDRyToLCkkQeHL33BYal6z2wpdWa0i4C9omeIbe8kLKWYbQYvOkQeML0zq1Zjaw
+HqOcoFJVO4e9Ag0m3COnK5KRFBj+8buF7a2h7rFMRVghLV5Z86Ed8leynxgBBVeLW4iUkMNpvAh
SrOxk1ZXSF7Z6e50RHe1gf5pZGuwz/jxAZLC6Zq+FzFu/PA0/L/HPrAKTtHEStuF0H+mjy4tiDS+
ILA2JHTNQGzKQsy8GPvBaIdZIue8Lpfjabtnnl3S5M5U4PzHEL+fdif1LqrAmYFygtPLXfFCE3SW
hry8/3lnwmCseGE5ejuOkpOYNJTae0N4YeurHwD9EsGZNOsxBZFzAUsjFJRQz4xbjIpdukAW9pfn
5baS05zeBGKHDlNnAj3UUw2N01g3GJ+QXbxFjCVl8JK6ECfT9g4Wb0jDJfd6mxQQHpsYVdnB12IM
y1cmEyC9ETE/0krvfndiKI8B/bh/2qKn4eQxrcc3SqbfRvIcYqkTqyaD8AisbslpdgEYojNHa3k7
yAInl0xJakRYz7tV+jdFNgy8NNx8YQ0nuuEfJMAkSlw0V4r1XTCRurIHjKiwCNczVkX98oEoGDL5
A9RS4YvVDxlb5UloIrn7oHu8PBh+i2MdSlMa5Mce0CkFlqmyqtApdDqofhFGuVUxzoUG7qeuioxT
UGTiRKn3mPNO4vEz+kjiaOsz9C1pO3EwbN/fb+8GXJAg8Lg5sJ9h0+uZUOv32M2sEVBa7b4Ib8xV
GcdKLxkavDQoSNdTtMbLuEVZo8ift1iG9sYK8m+Bf3qrgZ3N9gCVeIH7Ib6wbrdUAxeVntsD+Byt
UnEe+ONVX+GfgrOuKG0AyE0x8xE9QEht0FES0zua7J48MeOwFd1teHYzDEPTkFXecFQFHIBuep13
+ag1Lh5LFQJGaODSfelSjocQOgncQZZrAPAKIKbT78mUcJyAGTaoVsQPkL6eLNnYQ7S4teKBWCTV
ghNjRK1K4yFTMRuuMmn4H/BaWL1miCkCjUCfk3NoK+xGY85ThQ7t/F3Xt0fBfQekFTkVT0AEEjY5
hOUExQuFZyZUO08WhQh9Nmr1OunitOjC+UM7cE8LFK6ILYU69ObN9EmWEEyACNhkFnBGWLdkDbeK
OdRRm6kI+G5CGE8purtrsu92vIUnITpPyDbi0lsWnZXHl062efNrYGX1bzjsaf/ZUykYFhRj6lYt
xlHuAsbBhHmFnz48X7VTKwXW1Tlpn4TLo0/fEwiScXz24g0Hgdc+/YBupx/goKWySj/KdDwWjL6M
eg5YHvTsNHf9zzfVjaaBN1X7w8eVndrzbLyzdZx7lLjfOwpJ5DGmxZ+JXoGTBJHDYQ2H8p9s1SsY
fWFWheHo+0jB2+iNhS0gOEjzFCxBmc8IxqblMy2RTkI2/24OdGaUOsST262XDEQCPewjNyOi3TJo
Og9mRycqvhmZO2hOHo6BMFQJiXKvl7P+N3Tmh1RRls7P6FYY/OSK8oOxptR1QrqAluD4nKH0GRKK
NsXUKZtlL3ydjAeVSZ9DT+4JNtMTzS/HmdlXkWlCJ1V9/dALeDijYmIZD6kLj6xhMKuJ8nRINVnp
3k4SSrftCmrXqhmwhZEJihahou6tbvYUjvdIxCYvBGKX2ljX3Jkgvb0yKqqgmS1ob9OSd2p2iiA1
/S1v4bRcFAC/GbQBtSP7OO6I5yqRugoqLSRpxmRvS8pdtDwIHlUgLPTe4avXsI1h0o4oCqprIjsi
7GdV8CznNjblbDNEUdVIdcyLC734pj0WGlxNB5Z2AiEKZrxSyMaYTqFmnnfvYLujSmVF6e4xXd8o
nBKUaVXF/7kdWUEaGcEIKC0mS4+xt5LHSHm1Lqf68NGPSTXArbGwAO1ZHHOstETBMzULHUsqmxtn
kIYF41qu7ZlG/AdBLMFk6sB5VWOYBTPJ/ErH7ZiRlgQElwMLjmzEyNaOnm5rhn6BLT0cknKJNn++
YwlUQXEoKlO2LtAmBJ/UPc6XvxpcY6LBksU++BIT/qREwUtRsLaYAdVgJbzDaymwjxUJ/6l6DKxL
BfpR9+pDfj0YRQYsKS+qGoa1wJDolRDYuvMIIZbb6c7FNg5ppD0ewMFy70qFAvXzsS7Vx6n1X/ul
Ws5biR3B5s25RSONY+ChN1qZ8llbkbNE4jZPCB8ZpLJgwKmH/ju0DMSDYHpJO+iQPbd4WA5UtQo5
C/8fvh5F0Xksba7UQVrPDHJlbzL69eqlAImdF9H+Nz0wGXYu96xxDQ6QhERnC2wetNR7b+w/R/Ta
4XRY1b2EJUvT1p/j/TGVKhNk8JNoyln7LLksST3DdmYjwIjCcgPc29uQDeg4ycTGxd7rygeuWnuA
2hyG4yqcWLBqgBht5AAFhcI3ITrHNPIQBFQ9K33KcTRDf3HmF7997kP6QaM8GXATyKe3i1Hy6wix
yyAu0mUaMc5n++jcNslqDhWmm7gEI0C1PwqNoVlqq4EfZCNdnrAXYT2hL7opW5au+Ff5uWgoYqQo
1cxDHVoBI9JqWManBIogNDaoMxKh6Rp9ZCWAD7JpYeenV+OXYIZsbGd1uaSO8UuHZfhMKg8uOtFE
aJrub7+Qao7h2m4K6l7ytDqJEz6iGGeaTN48aJFBjbmNTRUEoZXZB/odZtFoG/dmfKex494Hy1A8
xLn/zv1T02oCej2KbFUj7s95FrKJwiozChjzQlEA/n7wci0wKNCr0Uuw3Dbkl5YN/BrRXTz2m9VV
csQfaDWU/C6AXXM3jl8KGoDCkoM/qKazkYal6QjFoO2/s5qdJm+kpZeW/edCMyoyqrzmg41aDwX7
6Gdkz834uaiQOCYvwP6pfdTA5rLAO5CvM1ivANpxQM9uAksS1IQNIz3Ah54N4JEFRTYhu7n8Hmml
A9egBer6L+PiZnQvon2fw6VYX1a4hopqMVQSLyTgETGFRqBq53oQOWA1JNsnvBvjE8RXmBysINuA
z01eIjhPF6mIFOm8O7x/rkc4yivZFZcMTMYowDXW2HQts55wQOiPcxIkxu0TxFGrpNODdlFTsg6b
BhqmQ66vSkY34NVnAIiAJekRGMBO/m0lX5n4jATZkurAN9AnlRyHqFplLjiKmeB6wb+kds/BwOL7
kpl2n2VHqkmK+9WR8jFfWnhzw/Uo8LCihE0kiZGQEwktr23pIRaHbPVo3SDUhxZ8sse/3M8nHMeS
co6Vt8TcYEl8+wWnwG8bb3HVHW4UtceQ9V87DQ9U4P5Gbny9rESlg6OD+jyAASYtHHWRrodObchC
WvRu0FVQlOdpceftLAHqSG6fQ/M3D1TiN2fuG82lWhfwo8BgkEWGui+sHo6kMoTo4zLwrtc7jOYb
7LJkbTXPBW0UjdEFmTUfxNvcQ58PNLNG0Nv12Djhr/5FsGYSP1B+STLnZJv6kfJwmVLkEBS3omh8
C26Vjk8NB2BxoXZlE4nHAsxbrlNaXrdpJn2NFfsLbSBfOlDA0OSJQocwTAX0OXn0/Vfcdw9allMP
im/ZYmkpP3qu/iCx/lGl6iy0bxI6kyv9Pr083q88k59VciUglYgK72yOxFm6stQXLX9t69y4oca4
s2D1ApgDF4U2f5J2W3bSkL3Ph4IQL4lt1UAwGW+2XCK44GGDg/a+8POIqMol2i5aopnqg+7LGbYX
gA/gNyQ0U4wpwc0L0RlyD8KQoBNiN7jQiFbOooMB35UiS1ErKGagga/pfCAE0KJm+FIgO/P2JfBL
eyzXxJQOY2GuOzsEXV0gGoontaGGnpZ9yheJONOAcT/BTYLHt5ub77UuSuM9/C3gZu8ELL2aTSZw
0wRUCLfaI0GMMfW2FiL1CzG2IUqtOBMPBat7qgbKAIFCWu7S+jNmMozOoeQqgZN64GJegGMcYXD2
VLQZd2mpiMj57OhhOnSsANyrUVWmP2Pmme15mGBXlVO0URPy9TizHgbwkOBwfB8qhI7xoHrsajqs
eIsWlIM3Cpoi2fYns9IHzWGn1MfJjFQuPSt+xtim6fH86GkI6uf7AuqmokEI2hCQtTFtHJl7Wt7I
Xn1pgo5WWEDIMb4g/esDOivIEo2kui2AgiMPxn7OEFfiMNEzMoCJ8t+6tARe+5hohtVAdFpKUodD
GVsAYM2iCvNuCDdQQsfkJWJlCzp95lZ9e7PFTlAa2befj8TeLDJ21SmmoKkDIODXYLitYJO9ranB
uWcTXv/b3wLHe/z5fq7ctZKNvLQ1w2UdWiFeukkjhbym2rXyZTZY/ujec5HVvkHyRLRuUBd3gt6w
8fHIyJc9cU0Yr68czPgIQHSwsNgmRq9cGzLsxU/eo6r4WD9IgP+VR1BAcvhhWLXxWm+Jx28rVH4m
flmr6mTEQo3MOBVCXsIXTm4uIh6VAzkYZOD+0G3avhwfiMX04AurXoZxaK+4SIX3MSd2RfcLzWga
GlTaKLy5Tw0M6QK9yOLMqrQHC66L2WwQ/rOOEZnlR/w+PY+AooMm6YvsDDWt5CUSKPFnAy6XXlFt
kGGX7okBvHfV+JUl90wNjnv0syJNDgDX3TiMMb8VR9DlA7TcnkwTKvHRPQ09lYsnJyzd3iS6qwVn
2ewNO6hNMSXfpvwCCWOiavm5sywfzP2ekS3kzERvOaepv0SX4Dv1OppgD92bFrItczuDRp32fqwM
Smj0riUH5506Bs8fjx5RZqLia4a460iz2zKswrXFSyCWccscNbJEnRorJndBCQTk+8coHqoWSn7H
0SZEOsrj6TD6hCCwi8vn362dw9JCSpF5YtLEQLsX6Hk3qcuzUkTrwk6ajgBJLafoYZ6AR/z6Q0us
FtZecfKUWnGf9X/6QUfogYLcbw3tsrFr4YXsMUN+y07/wvUsAPyCeEPZCAiNFmXBUjvuloafiug3
7t6n3v9WgKq+CwtBO/MKVN954FwhZ54Ile7S2cyQPMlirV+xwaKhQCJFbJ+orYGRxBXuJvrbBk6i
C3c55TeFAnRZRLyRvf7XW7jfZPpLNJgU7cdUjmX4e7N5vR2SYLXUHZ3p0FZarr828ves9iq3NCpN
v0t/PTDwXvL9W9MFnFMy/E0g+iAstEGkD/DrFT2z21DOvCTdLyxxZlUlXlHRhGuBvP9vNPFJI3nG
HsyWNTil5klMaR4aBANbOpPe9Q6qrC8f3JIDsecfCgLEr2h2EWb0/qQQy6ZqvobpKMNvX4C9BCB+
nihMnNk8yt8VH5m0UOrhcXFowXm3EWyuG9Nu3r3KLzbgJHQe/QadzW9IWZgqpsfOLvDN8rrIBQd9
my3bNV6CvVGy1MeKHluk1wrXaeHYzc4gdWyOvH0i4H10UYWYY7117Izfi7vg3+zT+XBnsy7ZW8wo
Suwc8gNtUMBRlCNIi7LlIPehgwNGGqb9zHKiyBJ45jlol46AxJSokQULr3Z2WALZ9ph0YDI63Bz4
R6zYqBsZSpSbwxJtDPZy8ngtQL80pW91DQasV2DqKFn/u5rmDTsI4NhxQl4g2MmER/YBfaWbhRFn
DqAKq3oLaF/hTdcghepRx4VFNzNryT+u8qHPPHIh67oBX2IBe20ZWtMx8XebsnziwPGyFJDadgcA
KtIB7EPwiFS8+6MhS2RKOb58W7fsgksgbiDb2yXUIBu6Jt62kZtWvtPRzlZ6aqJuy5GlUh/M7lAX
QNQ4U8Cx75ZBzOBAVTTI6/Q7Ib1Jo2DE05chF3EX0epqDGcZocV+n2TVzpVOTIktEbDkXMOkmhYy
WxXOuHVHBmDOCEdzdmEa3tKFwpdVY5rnepZmGWTxLJRI59SDeKD84wfuShQyO9vk4+ZrpuG7HuBg
VG1h7xG8dJ9PhMqYuD9/OmEMpBZBY30snuiMxFTHLdua24DfLBSOthJ2P2VnmQG1H647GZjogC03
LFlYFCN2N4jcgW/PuyUBz5MGQT/h6ZpWvXQXpe7KqTFaxbgy0f8nbZZithXy3gWjqf2UnnkIUChr
/sAJhObAeqgBYhLDk8ynMh/BwfeqHb4LHAQqNYuvr0XFXOdzeyYoRGKB9Ny9PiUe+DAbVXiAjAf2
L7U4nx1Em/zdBd8VaosSAW+Fw2a67t3KtyFZkhu4+OO92KoZcffFdKpUoG2Ffc2E3aZIuNn3G7ef
WUC5zCx8KyC5cobevbxQzfxWwqD+teORfQLhxZUmgPb78lvp4zFRyBIKl8D1B5tevFxi4Dul3amr
ZBTcKIu7TjtjqkyPoeoOjMjsSzrYM+4HG7H3IYOttpLdOFkX+1ES78SVTSK2MWqbsELdNAjWzBBO
vK1iRHQ7l6nE1qyhVimM4eKx3WKsPa1XzYdZu8R/IQoCVHlMvDh+VnAD8pg8Nk6i8zZ4WwyhMIFX
aaeIVKfJJ7ct9gtWhed81WMr1AmEiasPsKv0JBZ1t1rjxfDWb5OM8Ke9aCabqGAsQeYUNX7XgSw9
tqaesmzorlSYCzHXoy/D98svx35xFKtJvJQ9RXBsR/elUW9D4VwDUMQu0XdBFvHBbVIMP0ej+jw5
KglIi+FvU8LPQ9i++8lU33wUbsOlSE4WIrkJLXInZ1GffZr3cRGixG/fBT2Eb5ieT38hxf0mp0sR
hXlngPz1kJj85tR739Rzzdwgb/LCCZGDHS2KQgEwv3gN7elAnblL/CTencDP1yKetWSwSCDZPloC
rm3YHuvIkBYDXmYw8pcBEUelwDJfeKrl3Ohrh5pcF6vPKIqI+9VbkM0u1sCTJw/vnsqD2ogYVifV
ManescXmr53BMACJnQn9Iq9zbIbIzgyKkH7Oh/ZnZWbCdl9GAN36I2dzUcdFoPnDFWp8TbJY25L0
MNyEQSb5XEdXGtV+c8OaJww97Gsz91TH5VlavMQKY4bJj6HGsJvwUB1nVg/hplUe9sZKDgbjoqkl
5ossvSMM9LTwBWPFumrBnBGSQGXmz5i3TMNlJDvTzIA5gwKblaL6/0A8bjnBujCLhIVgaydowodl
XxvtHMqESbd9OGbf3YbwTLH69yGwcKq4YZsxKjZWvHfwysAdBngohxdDo+OI4Ke/m89ssAgsY8MR
DgQuomrqq8GA+9u6vhgb/FK8qPJHTo5gPPpipgQzlZ+dBljlyiu2d5qAhm7RsshhBf3RYqHgHT6b
9TA1lSsQ+puR4XqwuYfgtfPyL3Bfx7AD4u0dmu1NrSSG7Kx/Y1wTgJDDrmWjIcDGnnwGLSnax3AD
TtxFmNzO1TTvfvMsViOWV/b1oL3DERKNyxG9j0dGhFHRg/cIh1ziWZ/e/H7wsb1CTVjLfbI3fe8+
f3pCE1mT9qYlvbncVYoLgEKs5ipm/wzS26Xev7UwnaXkyGjVm1+ElVNS0VsZE6y8lig+bbbi5opm
/X5injMAXyJuLBgYnaAWgXqfgkOUnGzf2mGR6juT7qq9fecNqfo/moN1vVck440/AN+CuZBJyuGr
LnZM6A9E0J9YQQ4ZTJRtaZ1+vo069m4k3mCvCMW0OdZZa+tfvcsTQvz4YMUAVzHcALHViitHHKHw
SuHskY9R2HDCVhdLtDFXIgV9NaFn+yJARfnsIapeFCZx8Oe04Qnr/hOSY+ceH7UlfE60ctxES1+6
fiFtSYOnN9aDsbHfKSDSaijgRzOlWpYKwILiAT8b7Qd2nCz/RShgZmzPpCp1yJhKy1aIZUza2ohn
5TH9yg0bXa/UJgMTU9b6cZOluvqCa/XcrLmC6bXg0j8Vb+DO26SkfzwO12AnLs5apPRvSqruCkIt
77QlqklgXmYNyl9AwZF+nn6KlbYctUYupYY6VZ2VSHRn7yGptwfI7CtbLeRJ2Oet2Pc89yY9MNBy
qPjmrDRZZOSQbLUaXI9asJwqu68v0CfUe2kj3tq42FO2GJ11bYFAD1e0C6+IOzu47bLSttRFPeKf
L/C/aQZkHIpNWujJMNG89hic5xaoxph9dF1ywl/Udei4jR8HaK/7MGpmPW3HQDAKSu79+5eU2KRG
QdV5qomcSRiFCjqyZa6mwIHOp/qYKvZN32eaZ7Y6jF0hdpfdEga+06p/fgjWokipkTKK5d98do0V
suvFLoZ+MA48w4slh1cJoA3uLoVZ8iyvImEAbwUZUOp4Uzhw/Fi7pUxq4maYOFQ0Lc0rP3uQHZoU
TqefCsQlB934l2mQIaXVVVBD3yMuljptBi57813bTuOk3tsHs5Cn8FR4gppRPue4br+NffvDGm/s
do7Cc24ldhtxzfBQGOttGQ8lxex3bNOT/lPhKcSZIME69tEg1G3xjeJj7Evnbf9LE6kQz6yUsZAZ
+dMHVV57uyU/tgWJF8h4ZCoNX33aJGkMrjmcOP2SOi/QygbNyPUPttSNIX3Kz1SYsx5s20kM++ee
4RxQmxJw5YgBb1dHvfZZlRYDnFGRuWg2a6SmBbJMLjJR0jXskb0aohUHRXqrFqrs9CVqr7xr8JS1
ZsZ6nR3pbwKbqsOFnnEuGrorvYp2bgEjW45rSOQOL2L6Rps4sYVfeuiwtVXwMu45PL3XwM7DOw0n
cqVjYOP4BKslshEifJw1BxabHrXSDpmGpx5ERendwz3KRMasdJru7qWfUuatd66ZvqgyzeEVaaUQ
kKyf0CnIhzIsQqD3gr9uzsvfuq8W41obYWE74Ejo0iy7516aMcjuHFDhjfiMh1QqcuUwSuNs1VAr
FcCSanmWa5dRSfXEgjUh3tPyMB2zu5f4s0OKt2L4tLICTiXcdp8/Dvtv5xAYn2WqtHIz9XuRJaGE
MRVDHiqMc6jvQUV1qfqRfYQu0q5zBX9tTnn1xGKW0oXThSLgW3RCmkWvtyNm6yRSWuX6s0laGKqX
HfJ7jMOdoKOlWSQlWmxvp2CCK7kLuRJ35t+DMI8jS5fadboTZj87nfokpx9pF3eLU5Jxz9Iv/qtH
JfY3paAXsV4RVSrKxRGbxwiDj/gg1yBWZTYK14Ozz3CuVSUb4I/7IrGvmUfswj3BPuJepcA1BksL
5nqhD4sGraYNz+gCSBt+9mBMHowGpIREHP1VqJxmTXcPig0vyFsFDMxb3c4a9q0clnTU2vny91Rg
Hjtr4wpRCDO3IGV773wXThjXjLRMgZj/hKx+HYCUEGl9gvwG8OG8lqcrW1QI1nBU9xHsZY7NmQDw
NmmKtU2v/M12W8VOTEqZVLGE4xm56SJ0pPTmUJg61Lb/o0wsurxDqYPck3GjAdPSO1Ql+O2pRxUj
zoDKEPhNNfw2LAiRhiNHs/d19sk+4AG/WwjCzHe3QW9XLdaB/WFm3P5jlUmESRIO6f1RdFKI9Vjc
j2AVuU7FXQX/3ssCenO5/ycUsevkAAb+o8H17qQwLfc4PL+O3zLHeoKFwV7nYsul8H0I+oDy/XQo
P76oZQQ2Rk3PqAbraE8c7x+w/aJp652K7pIfB/3nraEx42FpPmTmgHkdU4ICb2VA1kmjLaLLKXrx
67Qtqre7mEBkcR8Cnr2Gi6uTh3/obi7tGEs1+TUZT7iDNU5glkOWa+p+URpzeb6sz5Dc8i69mgys
eEhruHBwWlY1rvSQGalQhiOLK95tLVkC4ZYK3+FtPBhT1RI9bbDG9prXWXGySf563qWXvfw4oGAg
1BW70BB78PekWQzy9cCuyC2KdFyko53rMHsOTx2HkZIHwPoPQqKVxhakTlyyneWiu/Z79WTJMEw3
8aJVqmTPUvqQtkxhZZoICrk3XA5Dk59ZzgOiaFambyMGI8fmgDE51CwnpD9vowljV07FWgfbDvMN
CDaxa9N3kKhy8wJl2aQp9yED2QnGUidEn9L9pAiGZaBxU2GQuWrArCs0kOT1VuBXHxfXRKn1BG1E
2wvLkX6H1RUiJQJR20B9+pNRiP1CO8Uc6BggtOKmTd1urD3wh6e7GO5jG0pJ6IdmDTjIxgEeqAtt
1F0HFaclEUoxoziuZSc2QWQAFitVPy2aZ3aCbiP1w0kHurMCcGf9RX7yBXUtRDm3OBTN3eVd/Z3h
nG0dRHuTUhShQF1yeSd8TN0nszY9YZiaN17baLl371uzVP18Ku5jjd/mZYoB2skDRy4JEw9543Mb
ogofI+DknGxaGLyniA5qKCWh0OUblolRL8I2mxx2FPvuttyn9/WqCL6kTMindQPYOz70Bxpt4sFo
DBjyNg46AbyE1Y1Pk72Jq/HiO4tEogoLcKiqS4/45v+QhWE3DQF67t6Pr5v1ROfKDkpTVzBZZLvH
aP8z6HeRVMco2rHoElgu5NXQdUQMjI7qagSXLS/CQBmVV3w7zu/3JvQnnv5Q2SylJjLVOqj514M6
NKbi5b7ih5YlHUOp22vHI4r7daA1orz65LMcbnaW0TkR6K6abx1f9iGaeR/hcs/0J/UfSdPu//+I
9zP0mfTY9RuYkQBR9tFrab6ceByWBsXA6IRubS+f/VtChfUQvhmychx2Xhjzyzh6H+Y+XSxKGAMR
Ssx+YqTWm/4dWSNoBluf7OsqcChEgOrIeozAhSSRhBbNjEBZ5Qzr7q6SX05jXM3x0BpLb1ZpfCjb
DXMe9njQjrQ/2MfMh8fhPM1hFQ89UoZ+o8k1fuEmF3Sxst2RrmH8rG6puX8QVT89j2Q0xxg07JW5
M8INBi8uW5wSLJge0jQCRbkCTPguDO5qP5nMmd74BB+AjIbP7gaowOS7vU7QUKSdabjKo+HYUcsk
dM3aOz5j2ydpCLfub0RUINRiPfeFKH+DfVE4gmjWQHmH6CVsIXYgTUuE/EogCS0cXWgYLCvpkVp1
TvIhYuR7zk8uf2lvxsSFtNWLxPGgEv5tbU96fQXss+Qc2ofQTTIOQPY34eE8nzjc1jFjxyWlTPWT
9YRskZGnTl6/LsH38w9Sh+rTlbkjwHEvoC/S/BHI+EdcWSVxvWAcV47TPgnVYKYk92Mc6VeXuFcO
mU33mvmzWnd9TnZhNB2mJpJDuqroT7VNJSkjQbCZ+ZeGQ8cys048IkMIY3RvMqo8LV3Al04Zglu9
D10xk0kUY8RjPzkQIWVeIiXLKQ2Bh8eIAPXQm9mInAcxHQZcGL2XLdEItoJLH8EhqWcpArPawHki
vmQBAHUQ0Gq4o7bTN32dQ8wMfRm7h2W303YeVi4o8eBcr7ubATXjN+dAcJj2AzMFDZjb1ptRH9uH
oJ4qwG4Bes6wlZ4pqPPHOzElyWonGiP8O3PlCGx2LsXuOXZwEMu+28W4hBEm3Pllgu84/epFEg61
QyANN7szfp/6YYLnioLL0S/aMks0xiuWtPS8mWB+5qEcSbLxoZQD36fGnsFlv70vqBtHKlM1Ndlq
LFSSpKqxKs2gC0UiX8l5pDmQuiqM5DRpvHKpKwjTq7FNPzXPD22H8t06BWXgNG4Rnmcmx7fxMawl
npCghsM5vTiqv0pLeEcrhsypqHKkHAVjBRGQqzTIxqnkwxM5kYfY2C3gei0xFPmsEdxFGDBDGkGs
xhVxtfz9DEUejDy0xW5ShI4zU/bdwH98z4QQSxoGMpeuCcVq4nkDzcSFgF7//19N+ExiBlQ6pVml
6o8k7kMdr09m8gtIxO3vTHkb/Nk3ISVsM6EgGNvz87AHBjE7QNcs9CiqwJV2Mp2qIGgRt8DyhFaf
qbUROBsb+ks6a3/IybUVzNurJSXLkZUIe6fpzQXnvjXvg9MBUYq2Q1t73Z3+fDZinjKK6tTYpOcp
/WXmJH1E8cmjJqDdVEHn38t5EGipwE9UP9xCE3ewF5/Qfji3uXHEImIQX/9ysbEVZY7tSrLriBRS
dL4lmABghCTADNDvcIa6h0TUrxVlGiAP1OsOnx8kOD16//CmQ8mo9w60fny4AJLIJjv78FUzvm0E
wSTFMwtlYXNmvE4sQT+Vum8WwNnC/YpTFgVqUZta+j79H8A8278K3dPqVnDuWBxg4JXdIpZUV/im
TOv9Tcet0X+w2gfmSDN1VIa41AmaZJkPTAyeE8BvsblVpp+juPIr4hCkGyHzr+NeB6XCegRPbJOQ
wqwzqnSOYShk3HViIInljyFeHQIygjv8V+k3nEMKhi0HNv2AXFAS4xAOJ6fwsHgmVvSe6ETYNWv9
Lc8rPOg0ahQQoLIQxM391wzkZ/1f+76mBu2yxiktWAY05Ccao1f+g1+a497E1uWumeV96QSTuwAE
bdq/3TSi35KS/MfJDxdV1cjDcXZBiV4IZ7WTbDjgcT7UdAwELh9r4IN5pnNliOyYbXuQc9j5QM6u
bbp0GDY7137AxUz9LghSf1igYDd0EogM+AYs71kv6ozE9Q/JanWiPOG5JFeF0dyRq1D/6ACg4yzh
xrqkpVwfTZG0DZcDdzkqGXquQYTTgKEf2bvgM6T0AIM2htjejn7ake6UiiKKOxo0PYGa5uAgUezK
fFkbXUsFf8yHXziNuSiKQEJTRDEXQOg4NsEjrrnfA176cKsvzeYq6k1j37K7HmYlRRV0VJ7/kSXh
dZSg5tPW+YuhnEvYXnJXHA79E3+qrRj7369nguz8/7p6KxLnNajPV7sfBlf2RGSMXs7frdAsEmJx
knwe6TXwCvR3eGgTAsu/KbC5cyzY6zgaDiPk0SezN/aD8/Dpgp50J2rH9lyf2Ws4fDEsSL/erp8h
9GtWTJgRrqFvoHNrsI6SIQOlpTBZ2ykPDH7mqHdXz0VaKrJ7a5vG8LWFdYb/EQBOzD5sKc1Iia6T
QhDt8P14KyRGDljbZvfQppHN7XNG18uDz0h9sV2DYSkS+sYyvE9YcGBbDYQbeZgi4D/2Bg61k6Eb
IDVjGI2umstxvnuPXh+TinV86PAElp2wLzZTQQVaMc/qnZSfGYet20MrWysVc6yFIBlgtumFL+EV
I2/6ZVYoddNUyvIKQ7Co/5SfJNrF5RRiYq6V+8X22xP1OHcs9+pFnlRVxiAdjD7i66Ptru2H0rhP
0nAi1KtnF/shijCajvLDn7XLtytY3Hn/S7fxyeB5hbcDhjGOzqB384YvDhWO0lKhO5fdWhEitoTG
8FLOl+w5rnAbfRdIShivv3dlGd0xljP0+zhnBC4WmfIBYamVS4o+VEEFYe6LArwUaRLjYyEeugzN
pLDYfpW/YvEs9XmeWiOOcxaGof/8ICCey1WcSqjOqZejDWiXyCzDG9+uJ4WwO/FhFsrg5DHpAEw0
bHi+O7u4ZH/XWE5UdMS7I5fNuiyKYxRbjWIDahArrpJHnFL7CUY6mbUxZYrrH0VuiXkASLFxuSSe
k1DjjRbdVKQhzj2bLREjgqaeP1lsRXNu3a+qa7Y4065kwRVwObYR5Y1ulGi2nEnC+D599Tk3UZ6Z
SAii6G5fuh58VfRARfCldYY4CP11kuO6mCUaK8wtlS55P8XehB8lgaFrjKG9e55KQg3zZvjz1W11
277+l73TkS5Io98vwweSrr6bpbH/lvzyC3Z0p5U8RbINfr1j+XX7J2TDQyU6wpoKtzzgq11M7CLr
dnG9Lx6KJMLSauontN7lxWg+ZQduY66LuZ7nWlQKYX0eAequAfm3tBWXpxWeuUXAyW9gwgLcrtdC
wOsmB/vWshr3qc8fiscF8fT3dcSrpcgIX0VnurwYtCeQURnQJVs8w+GAFooG4OUFSwJRf6lV8koQ
XX5uGVwPG0Fok/EorNCerEiyyKC/c1sZFLtX0zlinDI6+XDh3cua2KSTTXZIsjdqxM6OosC7VE0K
TWy3ITceZ1zFNT0G0SgLRfPNti8rkhibKIt0zGnAwMSv5Ql6rGTuos7456rsZsfcZVRzl3AKEtel
BkSkE+N2wDZS5h3BvNsSFNn7HhP69kEFo+2XjO4FgbEWA0sPOaa3J4wuwxezV4jO1whxoHmEG3oG
Knl5KW2mtzKlljCzl3utWrcRBJRAAIJLwee/DvWaU7ixz8nWy/IMxR0JBgRDjBpIVpcH2DtvO3jJ
2cVm0jJJgy/8S1n2ZOTQHRQ4vHerHFZH2s8t1+kmGTSmWaMdtYG4RrAyOFFdic7Okx60fOe0L6wV
R+aSqxAUVp71GlIQP6Mto6Mc/hOGK5KtFKjMZqHQQvyM50/lEKhuIKE0ABNJWbvHNKjw+3MBG4v5
oeP0wiFmdJ/F9BanOcQkW5EriKPwyQrSgrykWrlGUuPjQ6abMjlfCeolhNpUPkPv6/nL+EnPoUPs
aP/PNIvZRsSw+8EXtp7FB+7OL0mOEQXVa/jg3RD1Haex8LtsIMCA4erx0qKx/qNtFf2BF6EtkZVI
WrHs2KyqbWGDbylFXXps9thHg/HMWTveQ8P0S0yzqRk39/Wu1MYw5M7q2ZmcTb4lv6GbZl3NocFm
bgLAOc9tc0dkIaT8C/rafw23kTfbQXDPwV4n+AHqnsQzRDwUBe2i2ygXIWWUXMOA9VIF45urCUJM
MLrs+wQyapZuCT/wFmoQm0i82V6jhvYE8ovdqli0S8yAXTioQ9RUne0/cH+zb+oz10lKrllHfbVu
trEz2LYDWhv0GqX29nFspSdZIKQiqzAVOIAuCae0arTRVkYFZa8J7qypFN+giY92SKisFF/BL7VX
p7llG5giEIuImM/ik8rzZyFEeO3OwqdgvAoGP5+UjByI38lBMEWHx0WnHcbwMK9Pg3UtgHddaYGv
Suk93QPPZfmJoVk/1XNDKwz37sBTA4Sbusd/4WCssaqAEax5XXSICPe5OARhV4E+lXl7lBK2WRnK
EQNrQnyjDY8G3lbwzMov5i2nnC8I2nPBI3EIzikaO1kNr+8vBLTu00Ayy64NMEKr5hIXqlsHKiz8
6dSz4l6kARX9faSPwsGa+f/SltU2dM7DqBCQWDUClSCdxvvbQflx7YQhxxy5XxRNkFcL6Y2CRsaX
XNnkmbkDgH4n/41PMaXeLwfByAG6j3g2mMr4tsOAyAq7FxrZj45uMYxNjn6Bhqg6hG2/DzZ0anI5
caXGX38Ot+oD9HdHN9tHT2XQ3+UN+3/+K98tREIJLnSIIgnMdxiTwWv+hKJyC/H/9FIUX/5bBHyq
1WpJMykVSVFHvxmRtu82VxSUXMzu/Ok2h0hCqB8QgzlcYkCR2qK0C+xe+E0QyMHfeWgCLR3P6rUq
METxNmCnsyoA2L0SR3zYw61N0vAgf11PXzJ+HKsDucwkcJQKzhpM+3r/SAy3B+Mp7Dp0XhvyPs5I
e9oHyV8QVbaLUstaOjISq7svDq9ARzqA7A8tD/Q+xLRldnPqDKTGEY751FMk3+SS6tY3OzKg0BhI
Y4oqvXaEtW/ksSC6yvh2mefIB3n/cpR6Uw5fbc87LsGzHjQtLlaFu08Q/8FUgLCAZSUP0jaas1W+
eQWAzsb2tMoVvvmaC3ET4NKbzHaWny1sqgZrMgUS30vS7wWD8wBluw0X7WJ91ON5Y+6VV8WsxL8E
tdft5CI+bI0CYPYDEf87kgbwJ5xw8i0Yq9Lc3Z7QGlfx5y77mlVjaUcM/fsQKu6FdkD0H6ci2zRO
OK/k6apHAW9ePLIUnjG8W+a48p/mr3O87sr27tdJdRunBZxWiu3Qde1IrJekMd7e6k4OY0fh76pv
wDTzIvhjLo5dJE45Z6qIAXF92E5r8Spkt26E3egzCmbKfxlC75bzt8oIyYxDyH1Yw60QKQNNs+6Z
bBlkv1nrTfCLQOcw/dD5IqMq3EAKyl1/9joVBsPj5kEnWcm3Ox1bZfehTK0UyN2lIm0XhFHV7ulj
1eRaLpFJ2OKewBh3UoCoNYzoN4pOEdKtQ1Fd22wEigTkF9qoiEAryL6JdpyLa5rDV2HsROvwwBg2
B81ZpsH9US2IndMWJWAsgC6nNNo8g0E9jSZ66k0hexXvmRRg+lJgRcnV4NlEkBWzFWuoBc3Tmh6r
6cJLoh3r/D/+KFcwlsau3mhs2NvWeTuv1AVMbre567b4x4e9EsIx38lrkbK3585gWJmwZalokBPM
LY6m/F7KS9tlzLBAf5Wm0QNUs4C9v3RmjoeeFRJBlylCvmnZqDnuaAMNc0NviTJUzZxBQLwCP/1V
Y2Vp44wAIatzrpIV+UobvS2HAeMWrUa3/3a5dMKpDJtlpbwBlcb2qmnaFq5nOhzLCLv1S08CTZ8M
v6YCxlah/6oZYVuF22ouesNd9/9C6m0bFHdFdCr+HLnJtb8lWdzhnVxeioDw3H4MVPekLfRqfDbQ
wYoLhnj5McHVgU6lEM+37W+6qFuKZ2t1vHUFCK+Md/fBZZ/3qlmT+s51+mPTreg5OND7pHofYc6Y
9nPyh78ucThf4eL3dWzobkZHMGBL1el7LivyhxMJF5OSK/Ij4D+OYfBrh2Sna5ouGFYqhAdiP9kC
crtoz7M+DmzlE65YHmq7TKIYYCgRvK1+AXrbjiwxa9AJdvwi3jXICzg58QQH6QjwiRjX37spdvqc
0AsOQ/W4vsi7xeir+Hy4A7FZA1rZgSAna8LxkbuAS7e3fojzzHfAO4rNSAltNoP+tXoxDS2zeE3F
NWV/5JCSQJFJifZ9AmwaCWAJBf2YlXPwhMBPrXuESfVzXge7MjrytGDvoaWSU+VSACw6eX8hqXCK
CKk4z5UmzIi8sHiSnVrVj74lnK0pq97M/0hXirGuTCVnXP8wJnEZst6uRqRby/YlBm1wlSk5iAYh
9bCwhp7sAdxeUAO+MXCfRcKHgxqf4HLLt6AJObeJgqYOrS8/pAwt7eqrDEky9lI/eeXK3CTGOQoO
Cw243ar7jQLYVfWhghhIE+j6dPO4j9y/hpOs07U/LuwvhTNXCT0O8LLWeF24Qm3p8cvIWxJa9cob
SQDJ25yhxn0V0Ro5c15m5evu8OQqK6MStdsUIyH4YOx9tZ6OU64KUwCMDLQ2k/rMDeMDRi1aeZSs
7715kOrje5oXICW/brF+pQcs3CyY3XoU8wgtemsKV69y4x0Fqp97BFnd9q4rzWwoXkGxT4ZWtlK5
m86cNnjEm9nbVOyXsHg4W65aPyiuLaOegRLX8m63rEGWa4DjdjsXOjKNNVsJ36AIoXnF57BrUjms
Iw9TWTZwwLufPmqJX0gAw15gtYq/ooIx1gVJdbAYt4oJTT2mm3s3sqaPk6qbLIcZjF+Vor0Cpcu1
x7GlefXLtn2uDObbntvKGb1jAAbKycMutprRsdE9metKr+vRK2JhVlzorilKIBjt3A6EMyDxEFL0
63ph96aEWz2316uSVn6yHfcjf+FZxjh0Vdi6Uz7gNOl5EDAdYuPzi+UXQrJxA6c3GA7PQG9pHBBt
tGh7iPF3Qx/eGTvfy18eAppPXBn3/esRdjPzlKxSHEUYdTAi0lvEFBX8OWIeO5Ka6Tjb1L486IWP
+JgwCt54WE7J+7v6dD/65wm4A38GvOV73l4ATf35beqXkUxYRp9fFtlTBds4XyIXh7nsG4ukkOIU
7kcKa61n82r+2qPST3gBd0q8ARJzgSRk1OV/ubjTvMIjl2TiRJJEaex2SVa/IZJMqdAgdQr/fQcH
wdj4TYWdzMi4x+Jv3ssZDgFO7TezaHYWeLD/4wm6n+ZHGTCZB4+elSNznetHVy0kIlxVuBYMoKEo
1nN/QcqUMD4csM1Q3NpoJfoFZq3zXf9kLnzS+iyrrAeZnoaYdZLH3vVzhWQ8Llw1yWehjSTfDSim
vBm1eI3tRJ46b/OyhmLidYlZk6pw3LHzORVsQDRgZn2AbciqZ/nfZ6yo4KO6KneNX7gV6tF+x6/j
0MRPBwJqoBXO6LbPGyeAooinKOmp+betab+Bn+96Lh+Esr7Jax/ISY/j+LOzulq6+9wyOVJIS3RI
SzO+7VBQqAg16jkxQJ01iMGccc0F6bU4/Zn5mdtu4Mk6u49h7iL/mJpwlnVK9Gr9cCiRb6I30eiB
9s7oklO4z4dW/bgSCuCybDMmRfREgn51CWiCzj7Y1wEPLCWPdqnk/D/gm4Oj52ArRetbugkioL3Z
YFtsEXX+ZNgyztk9oUZ1yc/aTSFweWIgEfQJnyynt52caMbB8zGHuV6OOdrwy/zjoClcsV5DF1G/
eAHQihYYL0JTt4c2H5oFSohzKfMEs9FBzUa90Hih4/PtcfLKuIrTCXS5W8GC4+AEWPhKmRWcwCHE
IVfAICCImSpjk1+IrS+GZxS3srxbceIBP+y/zbweVC7+MDY/aKl9G97dUHlrYYKURTy09kUSQZPz
Zyi06imCgJOPajZ0/iQAeuQJ8aksdqmDJQdrYEa0AuNX8rgaqAtbqfCGjau7MUBLG7rhZgsQHDfh
caN3Yt4oPzotN2sjDNE75tSgxyyCqTqV1u7+KuLn9vhQkvT7Wsisln2q2OMQYaGZWbWzOiCDGp7X
q1hFo4JLfk4sdgDiorOazDH2TqRt02FQ1a21NUFl24LjyYqFoFcWeZdHW8lS9ztLqPhnt3AX+hLr
yi/Fhbq1eSMFzvBeMhSKjIk4Jw4kFQ+NK6BdODyGB7T9SPGGqSyQ1YniwcN8G//UmBr7iNPiNwqg
LLjcGq+tQMaHV6bvAgrxJ/Ggp8MumAd7tJcYsNK9biBLtOkglQTnUhhkd9HC27Mrsjtc5U37rdNE
mOgFinXO2gDnngvbU45i9Ul10AUEI0pijAZyi/quElH8iywMOFG6M8yLO1tfXZTsE+58f3kCRNz2
Ivs1hi6LpZMkGudh+hTNccdp0WjUjwDdwq7NsGlwnkZyIP3NqiIxN6ODw9sfIAAIY03dqDb1sx+u
PwknxZ8O1GwFF4kL3BhR6WrYYxmUAtTPdek8hRsEfOgSQENq88pAZGfcP5DYLTWvWwcSqfl/fVyX
nFeigRlb3//wp0o4wUrJwX+6Jh2JKi14yfNB4DYO29ZoG6b7jP1y54WE+RuFuiMTWHTsTZnfU1xR
wOJ2TcW+ctmNReISjFXTAmTkqddkajiv/tdpd7k+9kAqBv9XIky39yaO3hcSUusbc7/i3R6Bx4zs
Oomt1s5/7gP+j1VX008dwTQ/sa6r3o3+Bb7+k4J1BG5OlAg9P4fojIUkAPmkK+UUUy2HBwe65p/p
yR10rzgwKxKexcocbbUP3UAEeGy6Ii20+YA/QS/LkhWhmGpBEhEJmRJYfb5GyFRaykt2v3fymWPb
i45hreq1A8TbpXGioaPyot+BACBP92d6929Jyy4lmygL3d1KNgDPzmv9MICyv34GI05rfojwc1Yc
TM2y33ZTDgnpchOUC+kMyhfXzIb9pixPax5SglJIzLBvC88gWdrOrIxa9Y24ulcePJI6mjZ9sgFb
JLOHl3svaL0c5e3lKqbIqlZSpJJ5TGL1VJ5GKPgQ4wcDgGYcOaGP60Lg11ljsUr+iZDQFcR/BLHH
it9J7hMRbuqLbjSbPmFNIA9dxF2UHZaAfz9cr8gf4YVDhNu+Ivczy++vVYEQdSm/LwOqO8E3zX3j
upnBmQ+wlP3opomFaXWY3LDyAoUhgCTqHp3iKWf+5OrkCauAoXzhsAPJGekxbNTTAqRKUmX93emh
58enR93ioy6jXxdSQA0nbkyJ9TY8N0KYky5iLrGUaP0phbviJtXQBV4WywbEi8NKW9ZVtleAdJQb
XjZ2EXywZ1phZpu3XaNvzRocRS+gW1GJzt3LVOArefC67Hj55UkFXSXZiXrwfmWPXQrIPz8gey9V
TzcRG9L66Pra5Wl56Sct8GSIcAw6DuosGntoJ/jD1KRHlFa6OHUiIBzW+6e+v6AsPyeyHHJFt81M
WNA6QoBIdpxUPjbJhUzR/VIDlQ78j/XTJU/Dq/IdcZzrgMPtNoyr+Mn3xoWpkhcNXh0WZvXusvlV
7wcQ5TSTY4Tkcxz0wG2ZP1jPqQSJ+VxMtCCPkprN1TudcnoYIZI/gyqRU0neTt8qSSTt6tAbbmdO
8EQVOCCB8YcgQBWYD1xOqN/Qf83rDiTcbbD9nmtPFpc/ZiO8RUc4pbyr7JkH0lup+VXfqpRr69wQ
e3eO5f3JW7i7mVfdSnas+KgXBZiTufJ5Q6FOgdda1u1V0U8VogOfGej4FDsN5BsizLh3J3m0BY6h
JvSvF4eDcdChFwv3WB7tvZatlndwDoxbLg91y3XBpqpqS4zQBAxCqLRJrVu1c40G/ZhHpcmRsHxM
q575z0H+ibjSXeAQoyeIsscfs2dh4772158k13aMkrwZRpO4tiASYUL1z9vDUGJwS+rX4trO1lWp
O8dqP7veST2sam6Lrth2B2/kMG+peR9EZ+0wF6vWV1+/8A4vGb3YUWe6ZVPD4DAw6IgF8qcGyikS
E1hpGmvGO8DjUkbib1zImz5GAdHAch8MndC/2GV9p9cNLFjQyCwRXkus1HflAPOO3H+cVxpdZRyM
2RhstUYOrzZ4xyC7Rz98fK7i8WzPAHjN8Ffme/vlley3avuEs6DcLCtBhdnVWiWwkPKBbq+OePta
Hp40e8vRwcF5PDOU4r8Y2VxU+mE1s7psFTLKLKysrOqaK0iJVa8L2gHgauExDX8zZA7plUymJF4W
9DJrciS7PW/4BiS2LY/5NevbnYFPSEC1YCHvJNt7x7CxMhkWzM56okE6xMS/tixUF+PEmFAtlDIy
FnS9vs0TpmxHtu+axyEJCskkU5Xq3+bZVw4CmRSMOnR2WaaV5Fa6sPyLk2RB5j8v7dc3uH6vL5G3
V8nZhk0Y7fYLEEYBEGPmAm9jmTjAdu3dk4yLmkeqyUH3NOJbXo3gKqWeBvdCMbuHONBoLYWIn8O1
Ud5Fqu8bu9+2cRYQ4gW/uHb+KqLdtqnNFUw5svpuqyPLOUajUfzeQQA20Pk+YmeDb+GsS+AF3kUS
ppSy9V7hVXnCWkTV/m4j4nwfGqVwfPVeks04XEvBPcl+hoZawABuMQAdZpMyEVuC6IUVSqIyzC6X
fRdgajh/xYrUudx3h6i2YVx7rmdFB+k4G+UogMH3ELNKZpByUPpTgHx0HaK+lga59A3a8rbD1ktB
K+8AQKL95eBuM4XJi5F5C9kUUuzvCSvMMNjsYxrewO4cpz/qsv18db0fAXXYi+WwoFZdhh6HWQpf
vlMhRWTvH0gzkF2V73kS5LoskwXumUS9wa67HfoU64fgR4XoSnz66+WoJWVxcDwwpPfYpoae5o2A
5sOW9KNaeGTFhj0h4b3S47nbYldJoJZ3nlCbuYUeFZ0o0zuyk5xXeM0aOPEuPZbWl9aznqM0SSWm
bckuEmfjIGjamATZjAQAWMg4WGuF1uzZchbAMucmBKd3351+YlSlRbOkr5Cx+L6SXKFJGYmVG0SH
A/QPPRKwkaaOvEarg/n9CTPAkufWubvcvxFmVQ5J6zNqhQUbubmYBFwd7rhCuQYSIcPJOj+jWSx1
HxYVXewZBKiFXjUBtia/e+uXjIXfIV+n1kqAX+6iq4po+2px4nS7s1TGcmQJdWB3x6WLPStkny6o
MT1AQc2GkUqi0k4oayBw9s9axaAwzIDoPOjclqnxkwnpcev1Dia9Xz8eaXKo8vqN45nl4C/+v2n2
qNUspKi6Skm0JltEUqRTt1LnWCRCDoNPpMueg5PYRjBYuomZu3RQDJqafd7Z9F+9oIT2xzlew8ZZ
h6NdD8dvrbbInzq//XN61WuGnV5K9Pg7fvW+JPX8Fyt0Lurhi8ZtqccuLwSHC+98jSNZNFd4c6hU
3T3x9uQHO4KV0GcykEMLc8VSp6MUuwP61zv0y2TDxGcTWcZdFnG1lqN+WrQsKZiO+IIxZ080V1nc
4nw4UAaMgztzghlOWIvL67bMGDIrMKeISVnBZaELFX0PSzA9Nr6QRW/d7zeYiJK8IqNGkH4/m7M4
Io+lkiSNNL+pQnObBvUqNmsP0U0F8z0YE7bCmB4UgVrybfSCYnR/PGkkaYzkDvKnMM/Ie6x4i8Mx
Mwj5fQkpReIEWpL2ydrNUFncvtk2LydhiJxPKn5lqkwxq5wsvJHX6BMDfkxoJqLidaCeZRKbDCdP
xFKJ+EaBX5Mig+rG3muODFmYb8ruN9Cz4ue0f3yaPlMjhf2Ug0pdznpU1SXxWzI/XYHYaaBZhZin
dKJGs/k+foSTkIWWuNXZd8XQfIOyKeDLwbfwFpBclpCdOyKlJBD4zActH01tp9bOEsY/07Bm/K9D
qzhBWKeW/SyZ71oAtvS0nciHjBMlRqV9oJxYIlKhPCoWge0ZWJvOkq7gdO3UniiShe9hTmofmUZr
DTo9epqwLZ5FTYEZbtm35hywe85MGzmH2ZbrZbIvSHmGLt1TStpJfhkYEH7+KkQaEniguQBSAiDS
kCJjt4EYD41X91I6KXKexaAsv/kpSIfPFl1N+bexXSGpHwA2iex2yDSq6XJkBmT4GwHyvh3BBe40
swDjVThDIED4NfvSfx/MAS1nrY5N2LRYtK3jGZhioEtUejMiiJNhpG1/2oQxl1l+rpn3W+lNuPXl
ZtHpYO7sZgcDX21Dt+/3JKj7jkWizX7+BZYyeDjsxw89s5J71AnOMkaaSLqytBFpvhZ61jI+XVns
TgF5uhpQwpn06x8/LeT8mkeZNaxjBM9GUzO6WAKMB9Z3UEgG47K3x+V3v8ztXDj9jaJoQQ98auBM
MjTpJBR33v56wXs3R0s3h3s6NduQMLyC+DB8ScnBYDAgHk0JBoYsW0co0KdLU5I7lRyQlqTl5Lzw
odzaFFou1VI4pXUkVNrECGRxkPYLfRlsFVp+8rMOWF0GuOd59HkT3R+QuIme6+7PvJfTrWdPP1/w
X6wHTVeekAUEOWcr7U9mlauTBFvvkJxRy96eStOliu7wMytJYj35Y4gXczpoaWCMKSD/c5xouPMO
r4A/Ltc6QE10DM4xbiKk3Cw/aBvV8MLv6OHPlRlx5YcXFALtjzne5KG5sYKUauZaI1V4Cez693mE
I+hQnvIj2uEbYjqCt+uEO8e1rbfvCmK1LRUAaAhcSopgTvZYLl+2juqbymDlt9xpapNmS5rjVilI
B3/92N9BbKGVL1EezHwNGzy64mnggEKuPQMSr3w6y8cP1XnpaL1CegLu5cMqfFPFYbOHUr3xtJWK
eqU3JlnAnDV96WBPdMdxN4iJIYx/uCzH/LtATJsm/lJxJHJd7mSklv1xlQ5bHe9RgefFPI2q5xTu
gkvZPNvI/IGXvrGv9LFETJPLC2EGHbOKq4kOw2uYS/gl4HRfm3qHWV9+uf38NnlFw90koWtO8ltF
Ks4ZA97yo0qMK0gBlL5LSdhOlCH+azQozjRFYvgNgJV1Utt+wNubnrf+GmhlIcPKC7io53zasGAI
snhbUjaJQd9kViDnw9xDjFvUgXWWHxC7AU/NjDfr2Gtvb97K7lkyI+N5ciJFI37mUfcxS5sP/YMP
nXRml7fcWzFO4dMfK7m+0BicRBwhE1j19bjDaAXPORTmVJpiHWyIQrehNpLR6pR5WOhEaAfrDuWT
5/xMDsHuJbhgbUYQwwtKAIHnM3Lptxc6kBv8Dvff5ZceKyQ+rxKcn2Hi3tGI2m4FHdcE8he/yJFh
XB+KFVCBpy/6M+k0VCVxxhrYvNOF0uJLTnefrTRogQXE0DrWEe3tD/xwkXcD+MAs9OR55C9hqoHT
giYeRX9fT0g7JlI9iQjvCtXGlrF448fLGRI5nKWBbNksVt55D4wjsQR9tLoWIkwg2iikIPBZIKgW
OqvaqwfbnRalQ5UkACDR0sIWp+NdtSdgBpYGz4zG0sdRxWPCsOVuewNYM6FhOtOBl2GUjz71pAfd
17Ne4tlRe2YDq2puxWiLsyNbubwQksni9aacB+wBdSEslV2nP3J6aEikSnSpYLU1ZFSvtz7uCHDR
rlUpSEUmDI58gRh+v29OHZbko8UPTr7tT7Ih+BP/wkO1lUqKGvMlR3ci4ZiKBEMxZhY0j499rvB1
8rIJMqKDDig8hiwh9aE5G2F38otQzV57UTzSkd3cvnWJ2ySXKhF4BGxkmV+1NfyWrgws+XVf4Pq8
4BC/sLtvrmy8lRaPJvjwQ1dfWtRLgfFGLnXFe4URR6NZ2sFGxFqBZoZEIo+rjxrDi0UUVwy6q3fR
9djbgLtEM0iJQmB+qEjVScUvzUWyGYeGA14DpNtTtSbLGdNn6G6gRFguX8VrgVaVTCIIjg0TGByF
gfArio5VGmmXZyphe48M+EKzTqRSW1Nj6Lo9iFnp5kN8yXxjiCRYysBvuENhpWhC89S491MUJ6d4
ZCxadcpPv7yq4RZPoYa3ajlhn/5T+IJKZo4m8mZ0qZB/gX4NmOwaOfaRZ8uJ6JrRoluUTbwtSNzP
Ov0d0kyI4G+ANphm5K99h95w3oJLkMeiwrifVMNfgz9+yp6Q1xSIt2F77Fn4l6eGMTLlXoFOFeSU
Kg1K00/Z2LQl5TVk21ESGqYo8ucTFBuxU7XynLIhpfHm0tgAEdKh2U5HxfuuIj3sd2idlKIeekSj
1eB8JlKWcIxhUMEp/URH3KnB6MPwed6eg8m8ly9EDDhNuUYoBbavRtMbPRypIMVLYVPGt6vTnqFy
p5pyLbc57amqM0o9Dy0aTOq3ND8RGK7lewPtkFpr4qjzEzdrqXV6ISy8J2hsV4DGiYIUbHRAXkvw
M4JHtWFQsA69ZM/aLTRa+4aWxK3kktik67juuue6PJr3HUopRTzhgr66J8Z318ZPbPcmPx7AphKv
Mu4DS+S7GBfl3wwohxnHYulnUi07msbl3YncXl7/dwBtIsU0JsGfQRZg+hTN9bzaOZ0uK1JbjK2Y
mm2NabmxdYPzIBNP87Wt9NNpcjTy9ga1gtRbohA/p9fbpBo/ZmADzXt2NkdlhHwoboIEpI4mamao
ExRVkjvXLyaiDkBmBmmzxA0Mz0LFBsrdjvWqSkqFubQfDEeolChWeulhYqRMOkrCAXZ+mrE8lmZN
k2sqZR8DLwHaYPYfh6zbGOO0clESnX4xzwZLA6rpVLdk9UYt2gXANORXJhKN07Dn08N7MqsOcGpw
D7ZL4puBwkIUpXxPZUbyVjJ43QBgZBqhwMCA8js7hjfCwbXKAFU9NQdn6tD7/YpbzcoPwMwKA5mc
mc8go2mGDV2yADh0sxeUOiEqsfanqd540GhANYeLa9JIor6xqEjCs1fy7Z7qtZaNeW3l1S5B8/ZT
BGHbfP2reeS79fJUZveWt2pNiLTNXVAU2Y1hRQnYyKdBK0cTprxV+hfUKBV4uhwqeVtuP+3ep+cO
9d54AuDvgAUUNX8EldvVRB+vnaiRZx7iWPgYKlP4h12Aa3oxoQALP4T8TuSwTSs97YRN5iMA9lc8
qIrSGCZlR7sXTc6/+8mXkGcGk6xegUjm2smMTn2eH/+vPkUyYNsvma93jmNApvYhJ303qHO0dZc1
pdkpdIhkpZ8zDmqZRpcmYUjzweBfOk0AD9EYGMd8p3rcROiO0Ln5h1IZjRsHiJFpmPGEfCTvqEae
5qWzUsxwQsO17sm63ZoP20lWZPPt74xw1pg4b9073rtqsrBq6uRKPubRdAtqQ4eBZxZcTuY6C94t
W2p4Q69pK9szm+c/cOLhNeckPNXeulDfGsF0ZqYAHNeiD2jiCBmh3BQmIH+IpSv1efBDAz3pTcA9
XEQR3S8jkdj2WoHH17e1y0XE/GPWfHP8wXrITvRKWr/bTuIphK0Y8UPgav939lZkT2pU5EvnnCPx
rDefLR5IKRWXahrP8j4jf0epjMj+Hehzlr5wlyRptxHp7f7G2aBLYbxQZ/g6TaZQP3lkQ66hYVo3
/rc4JxYCcL4h0FM+1nL7NJpwBxqYB21CbAjnq1BQHxQx391ttp07ijHwtLsXxbwbjGgJLiUYlLUU
0lzVpjdW0tilsT1XTmiMfN07mbUpoPbVXruHpRvgtCKsf785EjfOQyFCphU5CUpFxETxpdyakoGj
MvK/e+QEihEmIG4nMB+eV9feSYLvQXUYxxPcHsP90pUt3EKrfRy7LGpsBpiwPjdEWvm60uBv6E8z
PQBs8dSiWYXkXzCcoMR4L6xHuLWpTT+Wn0mXP0/OYYLLg0GfduHpMM0ZDqWBUeGqn3aW1873Mqsq
uycmHuxmDfZ2r8+1XpYF2etQ19c6DoFKk21EK4x7/qAPXNSZjXbArDbn9A1yxTe3RclBtxFzQvUp
Wu6XPEJIXHoBHDFG9HAP2CyOe+ii+e4dIESOqNistu5OVJnM7bW9qtBELJfiyOGCvuee4IbXGzbg
YFwkWBDQfRE0U0sizn5KGtfrPc99w1jRHf16uQ4dCOMbFEPgqNk3grRoDEAmFndCsRX7HedXHTXl
OvdKbY9ePIPVPX8PpNxXBhCm38FYz8sZBbVt++hOUprugKYwcisFaVG18iND3ZyyjQTKDcS3Jklj
Bq++AjvgX9xnobRQIe/8B+1ofE/kaUwnFKFgfJIOOdvf3HVw5/yLoyBp3/M1cpc5PXbQpvdsPqr3
OMYrzk2uYhRVR7tplDDGOmLmcUkZBAQhvLAJfnk7uYbnzDpyng/QDwvaKqgdoxtZrpXLmpcAaD2g
sXEiEgKCcW/HYEdYdbr4z4Vnaw+/55jkYy1k3SADwNz7aqKIUakSDXwmAaXH45L296gogeDfclMi
5QJiMkxFKwKhWOWy4aQ3d2rSG5U2oPK6gIYhefZAz4Oshm6nmI5gOY8J2jdEGEZ/awt8HiwhOyWL
clYDtyaMeqSDnDlbeJocg4dY31WfSf2UfrcytykKzA/BTI677BIHZX+LR/PWoGvZjVuHv+sL/SAx
6JKIEgTnNX3kdkqTLFEQRKa6/d9U0w168DHcm8EEsU4Hj7JEszlBpm0VvTWfn/lSMlkCWOlkgq4y
gvpFqeEhFLzhio2rURJd7uLBW1bFVeFr4vqaKChgOd7LydclsruAA4XlSwAR+1z46KK4nJKiSQf/
bF73oYjZPoNszyck+hVK278Sk98JNZ8PMvchx6Rv8eJl9kYn1OLXsBklrNAglIK9hnZ2i2ahPBYP
sKqUTymH+BdAoKLEAh7rwhfPRZR3SQNA2UmWf5I72tLK7Tj/SNbb3NOzdiApYAsb3fti/2VxYtLz
B/J1Rlg0fUkS0pA98nCkcN/duWgKktbGT1Y5NsDHbvu1vw5HdocXNIAXn2Z5d9tqNKEoP6rpaxGc
6hkMYzNgCeh+kB/lfvDpw4qKgCBc6wws1sKoXFxxoPli/1LkxLSuhrXtmsIAz/NjuHRubFnb6sYj
YuUt5lr1nMjUG7l9Pi0N+6j+mgNEWqfiEJ5Ep3uMCFuWHjjbDHnDLWZDZ4CzA9klEcxuqYX0jY9r
a1sU9zED8dcTP0V0a5lLELgw2ulW/MVLUuLSS1YVpFirUo00iPKMX6Yf0g3drXoWpoZZtV5+dH3g
z2DgbyJXHAvWsaQd8ojLqkWpI6KtgtFYEmE0sUaNSiEhcpj1TotNhrLcvbpaXUZnmCaBd8mqcWZB
PD3nwJ7wThxtVpAIXk6pQ3MSNrVIwYNwg42GQhcQTzfLrOCQEyDrET5h9jbdG2LblBlokL09RvcR
tlL5b40HFEpuzPYd5JzFlcpQ2i0CvIunzyecXwQMwxxz4vC7JqVNXlFqmsEbX6PHlEAAJdLea0LO
xPio+3lFCVLXKy1/7zLakDuawmBVt1QxvNCYSWZed5uBx+tUsNSUPG6ToEu9BPNtr/eh0CTd11CK
6fh5tUM53qKrTkQQJJ83GLX06qfHrAJ7KsaMQHI7K76sQ/xpO22zTcIIkyeKefaNOA/oNpQXsUD6
2KKv25sZYvSEdujrJ/+7DGdLlZjHVNyQwsLe3TkHO/Y9XvZrBFXF1dZSEOFIOWb2oWgkXBjy3i5v
tImK8fok3AAgA7aFKgfw8PPxqR+eCDor2+Q+TqolOAPOfDghcRz7nlQODYRmHm1BtFMXJQ2JyXcK
ZjWWXRgjgqUFDzgdRhmiB5HmcvTPA9QBKHqmYwKGEH0bcvtpLATysPE+qJzegdcrIPXHfeESahDw
SThT10Wn79AiDB2y4Lic7Y50FzoaoHwse4R1idZpvnsx0J0UnKYsikh8vJZ2+pHhZ4cWuVRa7Vr1
YGFSFRTVCiSfPGHkBFdzxO/TBHCI2pGa5aDk41vNbFQSkpuPOzcARWb9qByatAkQzOVDT77KqX4n
ujWpWSLmYOGgeVK8AcmEiWlceORxXaMJpu0190lF/i/75nSUiG8OnrtbbrID4tvHNE+nSGO5Ug0/
S4UiYR6PFFWJwh5LzAUQo+7NmIoLoUbfliSr6BB2IUO62KbshmQTyqTxUZEO1tabuKI2HXGhw+k5
ps1ZEfPH/dI00a7OYnDZsLLVFsyz1mzaE+BoB0uAUNPhNbf57k9Ktm130FkEHjOuBUUSK/IFKJBs
Pcl96k55qzgBnG4C0MdribiICUcqbQOQIh1D+nSDkqyWhUhhaoL2G1qFaGMPPVMzpGiFPtmSU8KE
DOCIFBRCYSiFCKwmTaB3jiq3D1hpk2Vg6XaEcks7IS+j2sFCJ8kB13vDypcXtmiVUQHBv4vHs41j
niRNBITamEhYhki8tcx/60WsKbgcgPIb7O+xUgRd+Oo8/NmjTsS3n0STuX7WPmyagVGq7tBhM/Ir
9PzzinUW3kWyzXmSs14l0fx7smlE2IVLGermQg3i8RO8S/nFMSJKP8j4wOfE4N1g8G2DMuz34H5p
cWF8Omspj9+4sBXbWTCxryadQ2P4UY/+jr5lYuInTe7KXWqHqqwMeQ6jk+aa3BPD+1UJhVgXzt+O
evL6R1nOtXFKoMI4m7TaBoEheCNeKgD6WymhpsijmuXITHGDMPuI9+EbyAhIP+kimRATR3JY5sXo
NirJLGW2UjBO3KEHq9pvmadHmCNLr8llpj488tJGaDRH7rbVO8Sdpyomk1/HJ6s+cpHTaKxB3VOC
QN/fkMoYgBbPwnRJoUryTAhGV6KYbYLfCwe5NTRGM9PU8m8R/dMsKDis8l9t50NUYVhJorls8tOk
VerrVcdil1eJrlLc8Z/XsHsZRoLXK8fRWiEWHEI3cxbFhvWoO6dfZ31PrBxv+dRFpFsgKjbsL0al
VmdNjKNG99ONdOI1qir5xOobUi1QDoqatS3w/88SAybow+uCJOmtgqUek0KCbYxuAyKnoGC0mrOg
/QYv0MuDZRIjniCVoGCt6V6Zjnq1Ieqw4QjRCRkzJ79rebvhbWRbNd9CgaapYXWZzhQ+jRCAL7vu
a8mGu1zlZ+GZ+SzVch38Jx+MFcphCTvdbzwmNu1nvN72a4yQbyf8pwTpN39cdRhKglgk1Bp5WPTK
678ofi1ucvW7pj20uYg//8nmE/fsvnWXkP9FdkcPoJSe5TeJq4drXUlLyB+sj4p5JisEZ5hCwHxI
rgSjmK4TvHnvtr7mtGrl718OJcG103ozWZoTKLbFglg18AICvAAHiE0oE1wIsR+Hj9IpL5DjN+M+
/OwcJJQR6mb2gayRbCo+ijf98Cyi9iDmn7gWEmSYXSAoEckpIYNazv19Htq5bk2FWSQV+Dbr0GV9
BNRS7p5/wAV+QOhiCO+pSlXbgTvJWxwNUjFKcJin5Uast0SwGGdSoqxh93B8yV/Q0QjOpQtBN2Ga
OqO0b0pvsJydJXWjPH63x4I1PBgfw2ls45Zlf2B/WoyNH4oOegjDMOiQAujEdR5er6jTsKbJEEGg
yeHl4s8fSFKL4jnR7hrvbHl7ZgFq/IrdaRa3AR+IGoKafCYwhVsOAS4cpLMpDHGlbkGHRzT8gVlz
M3yZc4hSrNnbYrDu9DRAAheNJgblmLSbWw6fohQIIUhclfJUkB9dm6/uFkgpQGTUWO4x28V85Lqr
I5iZM4u/auy39JaEyKPRkjLHSVDOGdZ5c4gW9HceS/BfKgmnjG84QV1s3e91E1xiCvZBGhTqXMf6
bxrqSBmiDFh007KxPpmgxop04hUhxik6KXAUcVtqKcRJPGtGJ/+tOGP+hpzb/7qfFylVuMPPK+U5
piwBduvcs8cYxR8qcweOcdwSdxAgXa8X7TaI4YepWbf6JqOjY8d1Yz5CzezkS1vbD2jwGHIYUTLS
VifNmdZZ2uRGR0s8znF2mctvqdGP67uOcTjvOem5E0CJlhbB4RB6CKLY73i71kWMI8foYzDf8uu7
Y7yikOh/ug0MdyJpgVsD1YGDY0kW+q+hvzeYMYGYmKbrKT3FTcDcuMkU2yu9+yiI+5iZNDWYCC1a
ep7wwRdi+XADgLhg2R19RglhfcRkjsNj1KDke25p/tXnNJ+JwYDpB+l9rUD/teISbllA+bgu5FnE
+Y1nejsipBsfk0ZRGhB0+kM/pjQxFjC4cw0yvdJMelnPuSssP5wdHesJd3eWeJ1xliwi2p+WWPMD
feXGduRILgrqy1MHqTEEKefxV2ijcuWWF+VkJnif6gHgVpOz6KpI9hnMSo21tvYbIrJm89ljsYtG
18vH9MNkuGPXZ+le5pN56C8rWh75/LYtezsNJ/evqLlPwodEl5yjr/AKWjZtxno6O8kW7h7IJDGK
MBqtue3Xj7fVjDY7F99ju658xZePc9r0kisLq2s/sGW72JhcCLYu+7vaE4yQGzwoReqqDRqzlctS
YceOQ0niCj0CPiFaYf+/ZeRSH+DD8q4JW0pFj9NbrzHn3ruq1MYm5FGG1SwKGup40sQALDe5v8ZK
pcthYhWV8kSqF85+KJ07OOsjP75yiEeJrLW1J0fz5cGWBiAVdwmH7RJWLr+jppTwodRiDr9F/q0z
yUpDnikw/mRknLXe0aze1WSLKB2EnvjffU0SB7x3mv0lI71ds1Um7nal5s+1pfGo23sETSS5oYmh
0TLVs0tbtZUoEjyjHDisl4TbGi6CiimWRX2T0ToK0HolIhWLxTCW3LYlKJWhA2NyMnOdG5f6GSb8
cwzKkLTduLg1HSMR3oZdiXRIsNkXsignT0yIJMuh9YwYRwI+MSiZa80yB8Z0G08zlyS55I1w4Od5
QjEKz4vbniFLiYg3oXhc010wOh5tbg/kkDDWTw2kQIwy39Wvii4sxS4nYZi4giYaAYaB5xFtm0NR
Usqer0wzSvzz+hDW1m8FJiyd1Qn3ZVhl07pilVyqRpJiiqPNjH7dimChPWlWmx4A4M1jw62R0MIY
WbMjws/tGXgEQCFmp72r2issEcCIYU9re1SIweaRd9fX2CYvt5X9BshRC0Bhs7m+rvi5WJs4N34B
+6UABe2SfEjffTKThr35YlRSDYPPNTaXNpxMGFyPx3Wc8xhivQ8eZ2ieaYIPMDpshZqEyfnnAuUf
ixeXIdOZw2d7o4p/UNCzcn94ACxEKKP6FJDeYedg4qQnifec5Ob1Dpe7efPHmo0IJuG1NDfM4cRy
16MdzwP0+nOc2c8o2QTsnIrIZ4wWkaOrUyzd+rpn7DwGdI2CsCIe2lRBcs+xzY/LLgavxHVmQpap
EB+abFvHT5hGO5CJYF5tA6d9qq7wktG3LSUDvNi7xZ+MEhlXuUXvALDM3h2V3ucvtREAABQq7pIK
uSIPaMqAqc8jEmVCwuqRgo81lme7WV/PmuoRz9jQjXpBLrkB8yTYHU+Pg5re9Yxsn34l/YXkZw44
ZvaPmPDMvcFywgkyE2tNw3CE0PxgYKsJdscKPQYluKAr5jfckbeUnj+w1f6eqGBnwFlITIZiiMfc
SshljfQX3g/aQUQbES8o5Jb01ofI3fMAY3JBvuORmXPoGYcvkxGYDGgrPq9kQ50XSSb4T+IvTR/N
35k6bsJa6+qE2bAQoV1uQUTICr9GhhANKZuzrpOsoiWzxjxm8Op7XosglPHtOB8SGUsw4GOajIWD
qZGm8GGsyszSi5Fp03dF6GAf200ECHAkolY6c8yJ3c5sodrMWCOT2Flw87BtyUwCHuHvZPWmHWLn
DNMolpsKDyMr1V7ObfU6HdAdiJl2zZ2paMY/593ID12inkjy5qT4QdjXbttEf+8IVfpevAQowA+h
Le47yaxiQq0vc6djlejJJOsTIKUsFJKqBgZ2GN66VsD15mxO2bwqqxBFLhQ83p1Av+TLV6q7Goso
n8m0u/LGN1y1U/AIh0IyeDhomc6HgVNjWw2i+LObev9ZSu+FD3AcwPZVsf5aQO78IBnh+c+5F0c/
jH9SZ9tFRs/wHnaLlQxZxc3oIOr5k1Mk0P9LJupncvdj5x58cAOPA64VbEA8tiA/UGEGEDlwmK6P
ifgyzfYhuPO/rvE+Mspr52u2dfP7VEJiXNaYMxrWrbSgz5NjoqDTb+6Cm6lKZrYya4tRhN45eGKj
1a9imjBKqHU+inbPk5LfQBtmD0Tlwfa/HczVWWMn+TrWc0LjOlPdBG/fFia3ZD7F1GO0l9EMiNqc
HyfFrBCVfGby121R7fnY79QiDbFaCM9/k3iBSahAPMUEkycTdQkc+pOG0i/uJhRV24S2cGuxbRCH
2TPGkGMrV3Ul2hH9D41151iHnPXw1qvx1GYGswlm3Xgc2Y9QKEbYEJns1jCkf++STWXca/5NK1t8
GpyDh+8DdnwZ8Pr3L5/nJPJxle3Il/CTC+o0QYdeZeX01Y76JVrsDJT6VyqZF7z6RrMCAXYr22oI
7ZKxU8rOXjgnt2KvbpDCUhrTJQuuY7mtO1ibMWLPrOX50HjLyRWCp70+SalOXbyYo6O9A/rdWDDg
+D1IHKOawghzzdFNjkhtL9nfpe5jbqAIdQeBtLww7UTqla9Dkz2bmGLRWcBrQV9w894i0MNwY91O
nRFz5CeNZ1QkkHhyUHAciwlqDPLo3kh4RC1YI8upaXQth2esvL8mDKW/cd9xtgo72ozEW9uj57P4
5j5GyDaCrFUqNAtzRLqYibXvPeUN9TM/4Uy2YKSUqqL+/DqCK2p4BjLZgcUvBIbKHP6bFoaTnk5W
YxCow6ugjiYuV3DuHBHnl0Y7W7KkUuCh6wbOv2gfBQvDJXhAx5z/Geez31Z+YKqdLWpT0/R2xBjU
fQ52BcCQtCAOld5qq4+/rIFYMfxZXxQCfVgxaIvhLDsvFRQwkWFlsj+2adMoQv8tizrGHtQH4Xiy
L6dLyHsnXydmFWuoia6mx8TMrxEwmjKBktlyMQwxo8t+tgP7sgPWKacO6OEvYigdAY5J+yIa9rt5
AaLDuUD4DX8nRrLN/HAJvHzcy/OgtG2JrIZWzmGDGQXIt6iskIHQGsONTRO32Tjy+hNfkPRH5zaC
Cb3F2IDC9itxRK9JsvVafaXDWLldj7U4ioV7pCtIHqY08Z5qMu8OE4l+3HWGhLvt3PIFytIirUVY
YPsHNAyr8y03AAnitoMtt93bBh3eNwqG7w7CPJqDNshQT2OJV/sLfoDJW70Jq4Y07o47PQEALxbB
ntdwZZB0pWqWB4kCIAU8s5k//tuQkv1Rj5VP4/lquWS5ShuMtsGT21BZAcExFAQSKxhMjxyuDkLd
2/EUpNFe1k6S7KUs6gAjfisi1WlrWEOJEahDIPvEt1i7PT1GJEzhr/YH8viAER2RgvZ08L6wMGFD
Sly9wrWnty/DJ0PpHLTT0DQDzAYh5ICfrO0gp8U3Do+FOkfpLoT227nfk16FNHBetVCcGqnlHUJm
TlSu+H5hQdnjRKgaFIPG2t6nWu5TrFXPn4dfzidioK5E7TjOzjFGEyXymJJG0aPkoKRkhOXfyk3m
NyXV5Kf2OM5LWXWUJkDz0QriG713R5+FondMOq0SuyvKg7zAtJbhsCEZlmK6EWrYpR3vSOEom8zI
yKKniBgW005Dp1p3BnexxZCKkUWx6dzVGuFblL8F7MWWeW5afJr+6sr1DoaGRAoZPCrki22GRX6O
AQ8lq5PHXTJcOLiesosp5iOu9sU9x0K/ZkSG58QKhGJiyxAzDTBeu4+I++jTXor7WnrLKhXVvWDF
/F/QUPiEpQp9boN0uN4CbYWNe1GI6D4GXYmJxF/AX0d4gBePU3ij4ZrY6CKFPBAj373ym0l3/KHj
Xfa200+ssOuD5YEioZEbKDRdOyKq/guJHIDe5KzuGh3cf/lg7hmerZEPix7QBMyuo7FGddrXQ9n9
77Lv7KPWdBh62INkUVMMMbKjRBjWDBAdR0xnU+y+Xc4hlkPOAE6QMQxkDkFftDKn+fieh3VrsjwR
ITPqP/zPTBpJNNGz389Jyya0nsv59BpTlBc1YKepbKfcvgP4ho3xEUGlPzvSW6kUD7ebz6yetNH+
ymBB/zGG8lnlP2ddPU+Z0TnYD4n7jTY6rz5RqAtrRgtsNV6aBlUSJHXJf8BNev/xTra12cmegwn1
ZCamijREPOWVjkDihuxwBDbRdiCYmpm3QWL4HjOfcjc6ZK9nRezhYWP+TCiAevOWNmbLNxs/2GFl
/H/GRC2OKQmC6iW/TogNiKx+uV7BxTw/JGB4lqLnRKuA3OOE/bWRze3I3Ay8k0PSvJgyfmNsFpiU
epl1SUP+nmFexyQsDWFKEKtNtbhGlIDSy4wpKDCaTQlWNL9dJFadYQtHoGYeTs+N+yeUynfOdoMl
2r6rYw2w8g2TuXnH0aGLVxv3gHbg7kPxWKUsYMPiCuV0tyevHYdyqZw08OKk2Py9tdPKUjpIFfLM
hwws8DFXVp1x31nCDit7pO0f16RZBMY+PMwzOKS8hY1hpJAOnNUw9AhlIyw7tpNflBT/tQMEa0mZ
6PUNUTwR04+De6ItqxV8Fl3rWk0BN7qwoQ7MB9wlOO3w5k8bU2Z8ITRsTnpT3i0hHcKX7zDexRTI
Tlb8I+vu7+5PMcROMnsar6nMvniZfjmRobVF8qHcxKy1yIT7hyYKVI/v9hZ7QS/FS54FX4AIzdIC
7mJT6tXEeLiSd0tTTUgxy7hN23XaSYLsk9AMOJ/Fm3RnM/O1urapyYH42s3ads0PVhV6mqdjt8ld
TZV9bV7ApKqx4SO5zfxeekOT98jS4+yC+6Q3p1i/mo/lxyCF1klCLj8HLYt26ixob/6BfNbJuAIX
vJ91lEcXPEFDhbJQKeX4rL33iKtW3T9VXQL+ikh2IVHMfBBfdd0cyKDIpDM/YjGSOHECxBiuyDFt
YSwKEOYFTKkHTbZ+VVn5N/pugM5t/gDmIAbgqWgxHiuAJ9M+A8bKBpP+uQ5SpSFIn7y56ATLk+2P
rGvU/ptRVDyXYVuE9gVOGpe+1dFdsB78Co+uvZiLJER5kj3BcbiEvCLzffd7ghY088LlqCBsofti
l9MA33OUb6KD3TZNEtYk8btdaNTDup5TTUK9thUZt9FEkk8nrqz4dB4Vj/Tr/2MahXv3aRzNp6Iy
3exEqisOAWzWr4umSGOznewWyhEB/3wcxD/YMlgkFjcTjAFRrj+6FF6uSB3qjKQ9wODtlwmEd9we
VNM+DGYH4Xv3RqWVjQgO7DPTEIasr5yzzgV80GeQ9yK6vWwUhOLM3wngvoNGF7Nzwo8ZiveuUOTx
QmYEEJNPfFMz36Q6glcNIciy8Rcl/wFKJ/pl9LbWMlZ0EBRq/U11AZSAyq2dyw4OIdriBpyNXCE3
2PA2g86UZiE/E16xLsEiBYk3g9OFQPgVIC4FR6vKFm8GWiXFy5YiNexPLIfR5KbLNOEGGhL/sdAY
zIf/5nmDnlpEnJ9nTj3/uZVh2iWi3y4E+mRdJP1SrxmkVsN39nPxZLbUJ/MIKr//CNGhp7aTPYeX
2uF59+z4h0XzehIP7AwWSWAsBDxXMmF1Mn4ag6nr7fd4sbTnh6/xbr4W16tly5LonFwrFAAP9vLn
Pq7LulPRUodn6hPzOu7okS7anmX+h9M/pY0wGkkEZ3EW8ycZLIjftXrgkTv1lNB7tgPi17+LZU/a
O6SJSnuxzUCAN3A2MJqtlSl32c62G2XF0rhH0H3HlzmnfTO8O7ahewwwk2z768tuhM2Ph+OCbnHD
pTzs+AutaJLDjYo183bGXwdCgcs9Ul1iSOZBx+0i8/pkizwxol5XRP6cvlRPBrzsGke1sZYWlOxy
SsXjZuUa6Ej2J454uGfWNUuyax1hcdfOGDWY4AVIdJax41olKy2QoSt2vLYuuDJ3WKV27rlqQJNp
FBxgCkrS9OZwQc/vC3tltcujNArmllYbTBlPPkMx/y1ZL5VeKP2dBj1e54fQdtUW0NrRksmhVLw6
ijcUq1t1FgUKSLb/AAkxMgyNnjsAgafESdIMvODFRvlHzcPpPKWgSBzFTPkM6gxTBUFHQVwgGuNa
8aIRHxO5hee4Xm/u+3mTxJaoagjigKn13IJrzURScVmvhYcC65KfVAKZlxmrH3ZwdjTN+cYyHBtb
LoYB19Rg8vKMHLMPMyWJ3haE3eCoQcwtdSRbqr3WkPxd5gg4gDWT7TxYw0g3lmr9Fyq5cLbKvYUU
iFEEmqc0xRGxMsR10fZka8Ar612UEgc4JA+QkkesrnLF5lBZyzxZTDkLpNDebjjY0kmVLJ4lMj8R
tUJSLX6qF07SvHoSsplTJ8bSNZCEtwYVFwWXOV9RH/hekWdLXCSQ+bJOhLkZQoioQng+vJouNORp
RBbXswd2SHpEL8MD1/fUXykZO8Sa9PLrGSsqIV9WBxqiYW0OZyRjVhphft6l8qc2Nvd6imVQC8hz
AH66j9/F1vXtj0SxlfFuczipKpc7BxmpLhGfQmp70j3yXrKm5lQxMWSxU0DsH/vkbIsHSQ+MMkhM
fCEzBAzgTws32sEu4zUxLXcKisQBA4yXA73C9jcC5muZiqumAZ0Bfhdw8Oan2Fn8QPFMzWzL4ROO
uV1j/aoyOiaKxjtGVHl7hcKXg42rwc83WZbKhJRbphgM4tpVrJT6lWPSHuBK50mYzzWvC1a+h1Qd
7pNUbqC6hGH6ShVc8yJ/Es/X1DS/CPNVANXrLtXw7m/E1lDXRWmUAgotria0OyCJospcRyDKZK8Q
Nt2zMZ5TI1Ftd1xLo9a+0f/mLxZnSg2+7shjnnvFWwT1nrn9IDP7ZwmA+MekUWkXeEEGWISuWJQu
Srnmk7ROaGbcpahlNe1w+YdOGwc6NtCCmDAmvawCVrTwhSJAVeUiEsgKlhaBqNNWJ3/iaRY+yAqO
gc1LN3kDHJ4YcLB8MsJ9ULiunfvJezxLGa76w79XpTa+GmYLyjxwi1Sluu58llxMSBc/6uRQ95fj
iC5fx/rsINLpf9XQbgLNb3OKIj6n7FpX+kPFGzbzJWmdPlqqUNF9cRmtw+D+gl2Lwwdajl4g5cc0
g4lzSm6VjutAI2k0wlgwHV7TWEpyLc/vkDJTiEyZ1DLF5lUjHOih65629663xX3kQsBXRMHvVTgS
sxf/3dRy+mfI/dfA68sHCuPbIPslp5mtqQ5NDDm7dXXb3kSZXDWfDTbDqXyzoRKYBlBg36stl3yR
YyDcyw7+SeHGPQZWtg7u9m3bx3MOZAPJsInlZfg76uBEc+VQkQjJHL9+k1Jv6vB+poL4s4iwqjq6
KObg882QG+nKrqI58P8WNJeTsImDmLHRULEdPMC/J3Y40lejJY63WP9jwEobA0t79g9nrIaehPu6
FiXcAzbudyxTL9m65Ajq1vM0ortEJSpkCzhydqCfrBxC0nPQGxLMo7XOw7XEwqFgK+0wSKS7JZFu
D04ezWemdo69HaVQsa7NO0VAKJR0o5hA8Cxwu729m6NPit173GPd+A/pKe8LP/Ab1NKVZqEZ8ta6
Ok8PPnTWlcPT5qmd3Hi0wSxP53xrLx/1zCgzPmG9yUhU3KOZAmF2sbtDZqTv0noX6dbOYoIV7vTq
twpr2sYwJyIJOUkaBpN4eYowuKfe0cuV2dG/oKy45rFndcmam/ynx/lwZW2mjNI5eLspFvFeK2I9
5QpMR66EA4X3hQK7EAeGXv249fihmROTLzeiFOBH6TMnlX4rwLlBBhCPWlmqZ1azbd1J4/E2GMpp
zfnWdKl6NzFk2y2rGRv7IcBfDsLjvOLi9eCfmyxhnYPdUV6O2BOrYfezA0mY3LRtAPeMdH/laLAo
6s3288RjtSarGjUqCfJmo7CYTanWZOCzO6si3gsrj3BNATq3QXicr/MIcJ8bO3A5zT5LQfNqoyoR
N5RJTWnXPRljbDwx8KFO/BcFkh+nazps8PLFvj+FT3q/SwW6LN6YfEPvu4XEc29seN8LzALwShGv
eiNdfz4hBIVJP+YgfLimwU64/H1eG2djfG7AhgU6+cFRROT3/DCkQOev0dLV+E7j6o/0i2OzBtBu
cNCSFRDmx2KQpisX/6yzbf/KF4aA/+kfib98hmeqKiVht6S2kUF/zjooQByNgbSCmuRp3ktCnfFK
En7VnUV8+LHkIKkzNwxD76/7rfe/VDdMmXUqevXB4oLQz+Cl0rCfGASttMdMzV9O90svYN8zxR9V
OGNLGl0TGplD3oO8iJQdfH52v2+Km2mQ6SwAPF1jqzxWf06ccnvzCHAAS7aZoljgJf4dJgu/cLHl
FJv5OzyJ1+tIm42TpUIZji7AAQgQ2cjsCqVAsRdSZor3/Gq352uufkTaGO9XaVAJqXPXZx6U/PCl
hYQT3lgGReH0HC0JMzi2IQUTTmQ2fkzWT0nQcMaTlmbssNze7umPzA1T+kAo7AjQB+IDrMNfQ3Nb
y5mgLQuZXkNXW8p9EU6CcPbDZzuhQ2T8kczSHohcogfszeSpqKeCgYXlYy53VhHcJzQIDjaT4Xlu
D7Wc78E/C9DPinRKIGOSFcorvi7Vk9NDsD5z2Tj83MIkLxPc716OjpjTYc7oyt4etwdFwsIJFBKT
O6i1ZUHQ8ixU4uFgX0ytyvZNdpgaSP3L2u0iLgvjzrc+H6xsI0Er1wvY545QckUu3bI5qegIK2Ml
g2k2B60xR3C3UDCGeR9uHORWx6czQ9fcwxr5+K1354Jm2idekwppiFcGvbBWPWLSa0LuW9wiZ6qT
MLMjbBkP5QWjORMgAAeF1TYRgIx7LkekzE32Cb8zshV2TvAsCVU1XINoCGI+BV5sB/p2Xnbvywoo
glFYA5+JpjodPRbqBdQWcY13KcavoMe+ycRy6jT2KarteePD3OSs5e0ztBUlGHxAOoGu4cHqevYO
vFrZAFXydSYoYpi9S2ji78hNehXpY6iL4/v5nUaTRk1nwgDwuUuY5qf+ofBfyxVQqID+9Smmp0Tq
yktEkCYdH/iKOpkxfKmbv+yXQyJFYJdMqfti9KYKluxLQa+mFL/98NwBcSijUT/xeFP+Wc4sW71X
UussjkB44mjiBBnobKvvwNAxkgnyjMCJRR8+o8sbqhCUfkf37lxzCvkdk/4o+ahb4xP6faA8MvrV
zcl9+HPQev2uYxTkRltjpu+thVcHQFDbNFZk5vGRnUJ50Hf5yZu/j4+tS4eLypF1znxu92kgR+Ku
f647jk8Mmq7rDpopuGr6Zb+0dHV+fleK7L4Y8PkzxbiitxyBgX8Om7woCi0uA0o6A3BbHhsV1iSW
f9ebTJDdjxidWJWZzK7P1qeNudifJJVwYDDC7BPFwBJ+dYkRwT0W1D+EJnl/a+qol3Oh/ZhVLr+d
nm5ylCttQfcUNXZCgF9EXffCixbLYEoe5APhWlOp4IiNSWVOtaxHrV/92yOtUNJA5c/4Kosds4Bo
h6plIiPIHdpVPzOO0BMA1ufhwMe28uwev3UI9Bj/lplMzWJvc7u3+RCpFgPhZpbtuG6Lzv+0p0ww
ifZxZYKyiTAb97pvde93DIpeKJitOsQThaxeh1prmEtea4+kOFe4IuAuhUZYUCEQjOmjOO3xrhHN
xrweIOOUFvF29kc1q+RXXJxBEqWEMvDHxYFPojDUVK9hqT0s+DKYAZ4MO5A7v3NJh5Q22QsUJuZO
D2xjADfnMTbQP6zdoxHC5HCBSh3bJJsGylV10sWvesLlviHNJkD/CqQQnlcriCMRs6ZQEcfcCPZO
S9qh1TJ2hbwABYYRUyU6x8UcJzP126ZwgmwN7wHUVWZ9NTIy/lpaKZ64Yh1mstGGujNtAfDkIbu2
EQyeJmlcOqVeZ63DQSw6T28R3V1Z7Xpbz2F+a6wkbQGyBvf8xcLDQ74ytPu3c3Ge5JIPd3Nj2V00
a/ul0EAFzR/uqplNTHUaYkJDfEOJ7vV+S0ULBPyLEQXLtI5pWdxJWlubmmAJBTmNrs3MOfH2u1uj
46gG6n09Gxq62h7umYgPQ9daKVAlvRfvR/OyakSnAVcb3lbfiEGOflOr19O+oru6B3VswtYxiSXf
48OvVj3p/hBjS7aAePkW2mlaPA4B1F1jx8gjAi20UKhcMiWYrNbmU3h3qZRbubqX7iaKELn5RIAT
lcbIHSdH2iMyjNPQh+hSDHslzOD68+jp7Sq9KDU/iQFuXcIHx8lw6kTtRWal9xh76BKwi3x9h86D
AINR86Ovu8E5JUabOfm1L61Dpm8ycWDq3zPbaJxaYVzbr7n1RAkpWDAElKn0doGb0JIloNljajpq
FC9ORoLLnISVlMwm4aAsansIR0HXH4Rp8tgwDkiXj+4xa1XH560wPB0yCMqKt04ORkvagXbaZur5
30OcSwoQqbOdEX6PPrSFEmgZaGLdJeHsg6QSKWbhuBwxAkCfuHFHkslMnTJCeT7Ip8Y6w8nWaI4V
qKTGeeU+MEk40eTl+p9RAETFQcX7s0P/UbH5pATVRZxErgmikN5Y7m0rXsfPyvkSo8lr3iRW1w95
dLrYwpeGD4gR2qx0sFgSpPalMtbrNGYObUWtwXIcKlo1Fy11xkhIuej8k8a4gLuGw8JFetcKLity
maNmJUfxcOWHpHL+f6xwG1ir7Jb+NjgXQBDFVeKvQ1Q8+496wPF/rn8FF8zvLUSDLPLURxEoVsgJ
DsmjMWB3xqFKexVYc+E4y8FZ+cUG4oVkeh8PDvg0UCs5RKSW1BQirWltdVCUdZLO6qduf6oSNx8C
Ou9gCRQLZ4XU4+xNVyPXOhC1SBfaFMBoQqlin587w+dvQH5dH2xpPjl8OIs/UN14xEDJMEC3v/R9
/oSbwW2PdnWaXWE+dXQ5irLp+k6KiBtIeCC0iwpeB8mt9FHhuR1P41pNE974Rtc5q7YQbno5oUyu
K8tkDl2jFcSUXN4ci+tSGv+hYwAim+7EnKCHwHBGTJi8Q/R+ByTuaHGsXaI68D0ARQtWYymkny0u
J/TgA01SMpqWDLchZkY5sZmfFQmdUpJBKodz3W/xiqHK5ME5+QaQVA7ChA5hMxXpkiRg4ZGf143h
dhTqoIixvGqDtjqWcODd0FEhGf/17/qzH3X47qhXVCfLcwnjA4pCoNdGkrlCYA2/3GkpfsVle7qC
Q45gT6ZMjZbsFnmpBxzATZmOxvr73o802BLFpX15xPvGReW7R9OQnDRjr6rr3RC/0k7C8/Oc24RK
yvUM7vVCHky/mwunETa0Nuhi3qXUJA6ACd6W3MdmdQMhw0IogfU+38JGVhA7lURcm1q9e4xtE+f2
eSbp+PylKPM16x2m7y2NNt8iNghWr7UoK1CuceCdXL4h5G0z83hw7SCEs0gnUxTqgeVqtq0WWy7X
BXUYiTRJ9lxHpR4rIAfz2BR/P5JWB1lF8C+WSyarwd1m4CedHtbqv3n/WHKZfABd3VAbdpVd2+Ki
oibh/OP26TpkQfFfca/CCEgVdAC+EAMC1gcFX3ZKk5A2uo6cPaZadzsVFZPd2Q6T0F2x9dID2eGW
HVpIsMzFVjtk4BPVg19Rpn6aoqR2X87WGBsWaC/tGUZ8qLWuuaH2Y3MotpHtIkg5ZHyWWbOhDyVe
3+BlqXKlMysBPv0l99CKwSxRGU110m4/m7PtGzuDmfp4RSdLqXo+IjV434WMaw16Xh2x6t6x+xO2
ov16KwbwHNroBhroUHad2YOnB0KxZemJ65iqWhceg1imAtwsV85Ifp3CuJkNiAZPyVQ9Xx/exrWh
7Ov3yngE+2SvCbSoPl3ieHtSBIgDrqq5P456fx7/AbbRNqNSGCFd4zMzaJ2NVwB5KEEa/MG6bIf6
PVFS423bItCUZRwyagxrA3ghzVjh5l3W5STQxEAC00e0MnCut6HcXfA4ktjCNFj9ns9FdRBt0XkI
Opj3ofNo2AhB1p4fZLgSHDT+76WmWtkW0yvqXhi27PdDcZxGvlS+Ooqx34BC1mgQWU47kUM8GgLu
bNuZaWdUKzpiHVtbocubupFbujF4M3vabx6Y39SQIYZs+LUnaFJSzLyw8kX4GmWfAk7v+8UhzSiJ
K6DEpxpgga1wH1VIRVti/Q/BzT2hcIRvyxdXb4wPf5vlMrQa1rfSgM5iSZyMGZhI1i+IDJ0Bu3nW
NC0l+rVP2BzDZo/3LxsQjU1+6arGpcSr80SeNLc7UJUwRPNdan1ilWDOUB33Uv2VkRRGBGMZb8S5
M0LXt5rsBl9w1AZ9TvA2HEJWw0X9byzOMNUPLV7y1sdErWZR7BTP9tyL26S1moaZm8/9nZov+VAG
qeaa5dUp8Dxe/cGLVSnuXSSYoJvGCdWYxgfFumCCLePU++gBlaeb0ttaJgmeXavOugUPmOt+kr/g
8+TGa7jsPCDi0gTbLcPHyOSoD14oPxZSxoV4LHu+nLBlbaqUhunXFmSuZ7JjaGyq24W+it52V3ab
RBvTMsjn9vVivacULQX4YvX4ukfTOET/crqGC2pGNWtLSSpAtBpcE07VdEfcRFpTtsZ0TpGHbk+L
MqI5x8o0PF54sOStRUe6VfI46D5ilM7H7RzUpuWDwLQl74SnFDJbAL0lJZDrDkypvHZw2ZFXTlrD
mpjc5Ri3TtN6L51mb2uGqvrB9CbYR0Mnf6zNZCYXmjVZWKpnDyShoS6g9fEe+zBArnwrU9CEP6Qo
329gatrhhhKs4PbOPk/gqyYWVQBP21ugQgP90oVGmPT7gLA1iYCNtJP2ayx/ezxT067/E++jR9KE
f+QLo6375jb42qJdPkcaOkXzKgfYTtX7nGQ4g89DkeudLaTB/O9QJq4KzI8997O/YkQWTr8/v5ZV
aBYA9yHh1Got6Ew/YN6B1ATLzAyCZa3vDW73gxdnumR7uGE3k+Ib/K95xRUkG5nsHhacOWD8XMRK
mn9aYnOJfVUzvoQ9beZlh5PikmnHklQWb/QX4oaIc/7mHHMPmfTiy/0AZw7JDOWE4I/p/I8+AAGo
+eqBYnXNeGNJ/56Kk+E3vpI6s1WXnCIfvKNjVg6uvJONFlYRRkHlLYgKDSVWqhTmzCvI6frWMuwn
gXMlDEW8THWK6/SZgS2wYr6w+in0g4zkdXLpKkfCnayeFv0WEjDgCecqksfxJ5FnzU8vbp6wEUc8
1u980b3qsXRBaHXqvJtDtMCPvRPKT1Y+9ZBP6wTUi3WNifmfEpxpj41QYjsoY+BGGN1ZaRItrgDX
ypC+h5DXPCuL8wXz/dP5u7Om9NxURQyeZ1oZ/q42UP74+T0BGCZCbcfgpNAnd3AIU620k/VJmTEI
q7b5KgRleoLI7psY7Az2KpS9ZArwm3IKgChDlO7ImlqyfieoamNWnaBTT9mmebgTLQOejk2EtwPb
v325kOnSit+CyzpygrlLjR5Khfl/jmUfeMqXXOYsqLQGk3vARIImV4Dsc3goUkMH/xutYjPuYDRM
/fVFIcZVbjkpXjaUN6LrWHW+NWNSwGbce3JlYBN7jpyMvaM9GGwsbWtvXkovXMv8J1euos4N2Thz
8Do75wOgCDGXEn/2omrtXkaPbtUFglSR94C54qVncn251kDpje8AaRD3QAud2hFu92v1wkufIuFY
xCS73V0O3MLne8UU/ZSJ1RacmGIwA3DBqIfkCHzKh2ZRMZTXEf+fkwtdTSUfFhW/agcQuIBBCuid
mDi5GfVKcurCO4rGCdkwhWYdEkfkEwctMtaeneRHZk6ABv0rclcApi2axNQL+Ia9IoeYmOJ2JPyD
r/2Yw4Ul3zQuNLCAV+cjU8Hz6J6lcJY5qVgU7bzCq7ZN3P/SA57ILWhX6XVhBXi8Ego9ESBnqsWj
rDWnDRoMspdXi1T7sckFOoxylEb1M0+ymWKA1bTFaNLQbx+8cjutdi2ynL7h1A7VDir+Ki3378r/
qCMKQtaMeHuvBa8Fzy7nYCgDzAjCdBs9m1a+HCzIDR+bkE8Q30WsURimuEjHy6mPtCnwiekDsBMp
gScxPzd11ERYJqNeoDfQXN4P32VG5yzGeWkgwaChQNeWxHfD6oTshFY2uj0tiJyPY4ER39UPIvcV
Ta0H1oGxxHJnx4yZaGfIEQ7eHRaNY7ieeU1U9IF+8a6vNRqGWPyrBy6d4FeQmnXFIPIHxEwD7fKX
SSItVUOSCHSQ4X8sf64ItOvbZ7phE4Uqi0+JqpQ2DkkDbtCeXEBaz/3ll8nd6/rvJ23TzabBAgop
OizMXSgLrfpCyDvQibsn6MDyKhejo0+wHu6L3dymlTIRxbKnRkGOc9ApB6sd0XtD+1WlTpurLbY6
RmyA2t6nCwq6m19vGhl0ktk6cy80j2wOunVbuPHI7inW3Wvha5FucCOHiUw7CqcVHFP1wi22DVbQ
Na3dY22R8JtwAkWzN16y3qZbFFHc+KulnxpiSxxkjWgoH+OsvBMtogEKjFQa6KapcJadj/z6p1pb
5grJ285k06AJMcFjmgciOU1qDxUruw+MYGiaR0WbTty/uUpRUEzLpSoPd/vyb81ukrtlhFS9TuI8
YZyej8LRWL1Uned4yzcehLbuRFAfx6BQGAFloCc28RKw3Ml7puzhW4cr53letvg7J1kKXJG8FVEd
pY70BgohLlKOgs91O01FuOezcR7HDr4In3F2BF72+LNavTGN6l9QJFaUF+DXBwftYiEMKQyZRmx1
K45mmIq3rxgx9jOlZDG6EfNfMftXxJOQsXm/edVRp+rsYUnnhPLMDfn1eAVCFFxNABuupAynlabI
VFyt3G+puUvhuUUG0+OskxJbO6ilDuP7ED8fq22fGRhjeIkhY0ndWbvMOiV7wo4h2cSfAo2EP9DT
UG9UVv7P4qkj3DOD5iBWSoja4ote1Tps/d3jBPkYzzag8dnmGpr3XBRtvTT/Ne2z04Co96J4i2yt
5ltByBizm0T/6bDB5+2fH4bylDPUL81uLvlgYrYfCwBIuC4xW8ceO1cyqlwSx/rnUG3ZeQUfgib6
koVW1vLmlur1scVKw606emioLxZ4C50WXUj4sNF/X37so2C2elwgBpVIQV/Dz1qNEyDRvqXn4XfO
HP6ravPZN4a2+XO0iXPpiOlTdc/LJSa18nc0z/B5MIFCzXuTlfxnA5Depdohy3G7kDrzk8kXGtvB
prnqEZpGyx7duyNmF6vSErbK+OODOiTi38gpc0UkTnIVJU3fVt5Ua/8cezmNJLwuMcvkp0XXsHQa
B+a5G+33mYf0jQ1VuqEqs+uiZBI3elUYhRbBsSo0GgkPwAUh9dxRRb0L82/YlMR+4J6NFJOLmad+
Wdv/1srao4PLHN2g5ihmcfvyi1YONvA7r+Yrp3uWqM4jqXVb2FAxz68ikVQCZrQJEP39m8LBryIU
ouHeIr+nVVq9/W++IxJS8nw/YtLutHkdlQZ0PzwF1aMAe+fi/ZrCNo1MeQCFL80jIhLsgQSIcTXz
gxQH/C+T2yRZp/gpNW8vWPQpIIcpafs38ahYe/5SBskUsCVKYkTNX7mJVZyPQazvT4G5oghUulg0
P3JaYcW6MiZWHNUwhlk5Ts4HD4ETAi/Hr/Pp+ryQKYgJZ+IyAyhCrsKefUAldsTeFyOT/Mpe+O5X
/p8ndTDUmwied1KIhOMklzHAHqfgralskvx9HBbEIEhBz/j5USYRXExR4h/Zd3ke4t35PG92IbK3
SMQ0VtJ1LlLXMxCtKVa4yqjQR54oVDdiao8YYwDNihmZk2MB2dksVfSw3vHRa/FOybr7iVYWuR6x
2geFt9vVIkqpPyOfMx84cE1HuNRCNFKBZTtgc25QbREk6PDEfEdk71HeG+EGxQANeC/yr9RnwGlz
/FarRuD/lz54E4jx+eprOabNI+zTvQ7YGuv1twJ8FoeOH1dMzt1fAwnmFC4FzoCMpo++wZ8N3jK3
BLyrj0bvcnIMdMfRjQhMPJ7zcdH/8S3FpQT8Pr3B0Gwg3WZVK47Ehk0kV9esJAAxU3E68T2qHQ+2
DWncpcM/qOGU9GjyUmHQw5KYCuEYSXwE74YtFiTCi+MqqoiMiJGKAIMErgdjiyEE2jZ87OJ63cB/
XErzSvyuwk7s/1LNwIDv5JmmmM49OhJ/U6MGRtyKVG1tIojizPgBhycfy//TO/vPJ30Im6MZgL39
b0Kwqlu9fMGbP9Vu/G9GvlzJR5suiHdSYav5bjShKkcVsBwz2F61H4GfnW6gnqwxYBUsQp4aGsi0
MfB0zHpoN91Bu7++nqtXbDKGtckOqD0D1gMKR2XBIq5fs4Ymy+EuKpZbzZ4ylZ37/VuzzALvUluW
XTNUtdIA0RZ4tcAuZ48/G9XGV3jrepaL2EId0Vw/J13/z4vXU02mtCegcX2kdPQHnizfYfKyVQlp
ipyfzjBpBcKKHPuk5caherS+1RaKtCQxS2+fs6wQhtbZBo3aDCvfKabE4U8Z4mH54oEre0CcmKWX
A0T8NJZbfW93A3Va9LH4Dof6dn5p7LL1o2qDQJmLTl2r83pZ1KCOCd5z5qws7Jc3Vu6EBxEFu2A9
YOK8rDvIss3WdRNR+/Rmn1RiFGXkqIdBlvExMwzIuHPzUcgN5JFwNBsWGbS8ZKfLIfsplhVTrBCm
DQQK2FvTTcdacgt0Cb1jrpY6eloLnv7ERWVhUKjoND0UOQIf4BfUSplmeJAJ2/4jEqcYVJjeYEzd
POFHmhIZQ6DY0S6eCBebUFSgN+0b4uA+WcnHPW2Nbkwi48z4Y6oS3xBUpVTw4rypMIr1Taxunp2T
ErrYd4/VINstSXYL68OyOaqjcMRb/pwaScmrc2ycAhOM27C0RjRLmurTqIz7r9lP0S2o5EK329BD
d/s9qqEcEoelbk5db7QRVVpPegnHMN0qTZMH/rvidxLN0oNHUtmjazS47Df35zODzB/+sPrEBz2R
eVy2CQI3a/7uKkNuDzjSATGriA/GeRaoYslYEoSjI0kxU3/uq12mKPcB9AG4EsE21dKmoKyPKMe9
6LLwdL+7pBsxvyueTNH8BwNxvCuEB9jpjyHpA78v7ULPueuXxUDoa2ikytNSx9GXZ5FYeb+JnonU
OpDLLGpUX5jKJPnleThlmf7hPD0m4y24LKUEz8/WO9x97YgeAB0OvVDI3FueTxlkN5MHrBsFyyfl
ld1XDKfAIwfviPk+l8czvQ40tQ4xhUNx59ixWP8pbBgLxam/HAR43GPYwFt3ZpxUkuhHqvPsS/Kj
4ULCLhkw8DbSSjwiiX4vOklXkLos0RzD3X4ViqD+rjvwtj1EUR9/qc2nHbFpdrwLye93Z9fuUKl9
0gH7aRhWhUJXmlkg2W7AGbE5HyKO+KggHC2Y0Tm1sxpKVU+0bvV64JrY8Rat8GSL7IL09La4W0OF
Ej4iv85zs33QSZQ53lLRX5euZJinyVcCxuRBfrVavlXW4oQvJqvOB18UDShXv1MF7YcF0wGDDxfR
KLRr8Oeahr/QCACRIVA4nKxjFMLg0FBmLsFhC1YNBUKUp+MCeN3Ufe8jBEAFto0g+RrWIICX98dV
EIFsUURLF6kldOlAkMumP6otPvmT4fpa9E6ctt6CyCMtY7/xQ9LpkLD+vHnDR7F7o4ZjrhNzDsqk
m2eF4RUyGRnwRfxIwTtiT9JGA/4oQQEDfue5DLs7OGnEww99ibiUKViZnFvRqH87LCvdLD+bfQxb
kmTxfKh7AtidwExxf1Gz6BCTyiI9kEw4eWMdLLg620Sni7D9HsOdWl+MMxHDCyHZRYvXr0D3d/9J
F0WeKSRz9GMWpj6EFB0SrVWWqt0x5n0Db8oTw17tp5KseC7dZYLnjq4TK6yiJxyx5aLZ1rsOKtbF
evKmCcsgmouz3i9VoCPHr+1+MQ8Rp3EQdDGQ5xSwNFXfzFTntsdCu2XntE27EoJq8/q4zzUfFZlv
FYNDdjlFZ92YacXWp9OiAOj9bccTQkq1wwFsj3wIQpd5GotWDEODo6cYCtXi8Lzi/gkGdXRIZckg
8ej0QQRlxrkmcjprGAHeN1c/yJ1xZR4ZVEzTCc42e8KvLjawTi4hcdn2MBLIMQdgpxcg+IygtKhi
KNStFoKrLIcGQwXaSyKG3TZPTeHWVb9DCgNyHRF3GbFPr3dTh+ttYVy4PHk60hf+jzNFOH011PwN
RSSty6mKamcAOHPCd6E+f+BhEHv9dHaIoz1EhPp381HC8q2hTYIHhOg50rG0+pdSCCDuMN1Ejfjt
TdFoW6fxYMpyB1QjSuaWZry58cKD5H+X/Zi9aTBtR5AySDvcnOy/7jN9DV1IrebljGLz98vzH2sO
4VJ6uhRjHA6D0MmX6O7pQcLHQ3MM3A9f4jK3Y1JNP1QU/Z1svhwEFr3sc2wnkLndzhED7FkboOEm
2XtIMEAdzJNdsrpkDcW+EK47VK5wUQwZ85wO9dPYyMYjONMV98KjKtKGjV3z7VW1zJM/kCwCjFDk
gD6utgljqfaTr74eiVI+VAMJeXWeZLQg+tiY0ROskQOp431Bxmk4TSo1ffznLF42dFOJjCZKy8dQ
9XsT91+sZacYSMV2LaqSnzHfD1SVDi9Sn4D6oZFZ+esN3YClsA+iPpwbH7hJhSH1BH2VeQolY27K
aEXSaUu4DVR5vK4yNK01hGefO92ghOVVkUmg7vX/+MrvtPhgJtS3vqi175Mfo5Cv8WH5WzRQdt+V
EGUV/BWqY7I+ClvwfEa+8qyU3m+NFsmYyu3CXRlF4sw0fuY7H8kRLwYi84t6Sx7L718Os2aXQaNM
+CXxNUMzUFjU5sb3BdZ+KqLnt8xltIopMDTigpgTLaF82kRd+0deH2VVJnCVO0KNa5iqnqlJnVD1
Ewb0NIMrFLVt5me/1038AntcM4Looxy9BXCgvCIRMiQIgta53guYaka6n5NeXr6gYgRPjD7YJsf1
iUfNZS1onjfsyefgenTSYWuArgVG5vHZMAI1HpdNiG/yJcH7v6NVj9IY4ZIykw0IkeR9HFxsqXBr
KGbr9xdpN7Dr8MI3Rg166Lza+/l5KUp3xEF+7nVTIWbYd8G/D3lHlRZmPwPt+1r5fGeYSpUux7AF
0bMb7docwQsSa8hwqfWGUdhgx1LuKKt17sUymWO2htYniL0NZIzZcYGXsP7xvhuj34ndit6c9Dti
QV7vj4akXfnrbpFaiMKe8PcVO+Vu2QKXlLdMw+Z4u8O3mISKe06LPVzs4juEhmh+DfWAOhrZv6GE
mumw6vOMDSLVTZhIA6du5QQnrNcQT8Aj0KnpNT0YRSipLHob+Wn6ghII/U0rQeGiagKPzTWocqcM
Bojs6ooggYa7k2qvWCdOEAmROuLpi3ROQN9jN04ClDeZu5w6odfHBqwLIIOpo8VUyz5dhzZHcq3b
mq5zv2yU4MVtV2pZ3ky4qXDuavxzMEEb8bE+H3+g56vF9Q+nM1E50xnAlsDTOxqGRPRC2HKQvICJ
z57chI3V9/Up8uzHuVYoFyPCVFPMmlZfHzqecs7hUpR68kyQqYkGlfhUPgX8K1ZBaUGHpPm5MBGQ
y3+4us41clLXFvBic23GqlZqw5v2xXPH3Vu21tX+I5TTavVun6/RfzhKtafhvK/0k2ujkLpf2HCI
IHr8ZmReHkU4I3z91oWp+51Im0gYNB4BPxs6diGjUADdEwRgjwahD3fCiefMg1hVZ6WLOQ7bZxfw
KAAeN0akHQxD4BoI6v7VBCSWozv6tndnKbcqYlLe1D6BbHbtrv1ueVc0xpTO+yrleMmfTSENdWxQ
Eik+44f2vrePby/Uvq3I4p61CV2gJwOmnL4WIpI27Qa2LHsSVsbD9AZCZpRWVREp3McEYDuWnOuf
BQSPRYW44ZasMr/boxLK+MYambUf+C/AxVX6GyTrXeG5VaNxE4/2DCiAF9QexxJ/b9ctArgg0sDw
KbCU8Oo69L43V1GdRiof65Dyjr//iIOpJHBluZQzDeMR0Kv3+hmNmb8NSOP/LH4JcYtAomGNEHYY
FA7FMyStwqHLONmx4CzbbG1UD15dMj+TIiyYnqNOEPe2tF5vhd8HKfAGgpvA5Si3eDch+2yxYyFb
yRvB57Za8VZMmQj34ubVt0dzFE52vfsSZywhXvKmSiI70bVeoAFzP/YFCWzvAzHQqyCK+PlyjLtG
oGfG5MllkD0Mf+3BaAcislmxbfgQtwTMxJsjW9CgyN0Gn9Hcf05WC35+UlNEVj33BCfywL81hF23
PAW9/vzMOkFb7y+IFmITwPY69BsP93pNzG2Cf97Ber69E/L0w1Swq1jhA6URXWP3iSXCyI04b0P9
zDhRM/UTZeOCDhS7gxc/WNKr31dQ+fmat1KvD7zVIzaU62ZyxuD3m4B1Cu3ILPToCP3ARZdqX/mk
c53mOQNj711FAiWxpcQv1gsd+e9wIGdtr3/WI/KtxAsx8hOoiBBpaS+rsLlRUcBRdO2hdJpPQ8bU
XO66JgWjBhtmmz8TtX90RqCXXgtUOwrVPQ7XDcsxRmH0fptz1/1tSdgqPAI46EYRI4oI+fnY6yAs
VypZAci2mphO4KdyLQVtGZXUoPh8o6VEH7O1aoQZc0fbvGxvZaWwpyGL8qQWIVgT0NAx/xg1dyqb
/pdcB8a2Z/yDzRMZ8OV/VKH2pEXu7XnPz5ymkL0WoTaY91JgbrFVngqxX7SA0+C7ElRU+3LfNN1C
BnPOoV5iyLYMN9OAsLHSfBujgfT49xYuSEuwmNY1ySayXYTZvUHBAyM9s0F6ycgk7CzzGtKJYN+I
vdsnC0NNUScmdymzLq8t7bwh8hmvmiawYohCRG3WU2gSSXGyKSaOqhkap6NlXZMPd3Nc2hWPoMSw
sUx7+lvNucj5/NCK6+7F2B/SGENAPI0DsRZ5nVAsvW6SzqgsZlqFJ1I4qp+JndtDR/y1ztS0KFP7
9Zkh+7hAbjbtztIpNuYNoN4ywi0GJAJeYIijbTq3w28YGkU6RrNQYf5vcJGp3ORNa8xf24X7u21U
zMlVX+227HN/sI8dIpZiFtP2MiT0n+XCFloAEsgBxH5jxF41nBGm/TdUspyUIBhvAcAMevoZWMb+
Yr/eknVGYsvOlw3ThrOKN+i0g6JnFSp56egXSTSQptBY70LKPhd7SDg0XOEdnxE6umEXpxlYsDFC
WQQpSjttllx76RTzPFOwB3QJnZY7ExRgayo6B2BXPC4F/3fycCEyHt03sTFK9W3ejiPJo5lKPBBo
HWT2BjoJ7zaMUvLkUs8NvsikcYqjhI7St7Xo2U+2BYE+gRzwzDVjlwkuXoXjeG3J/vCHuhTdzcSc
PFm5m/RRURhD3lMXAnv1m8/pWSuooXdcgrpPMCA37YImM+Fuf076tBPuBKSfXgRaEwWp0fzzFxPv
mgQc19ucvUVPgLDKxL6Chc81GnA8mhpqPfrVV2V8mCTt35w4UCjuIONHHvGDoVZvp04vZpWb0KCS
ZAAM05+GN6tXmPQyJFWwelSDcE6HyTY0HRR2ybG11gnRKMejM+Y2/YV70LFzVanXQJQf+LZZlqeO
XTyeabCjHSEGeE5Kmb60QQmyXywGVcGK134CZxjevQlKRrY1ImUmGo5rTAToZcUc308vy6ZoEwx2
IpEu0IiCLfyaJUlvzS/r5zfMTY/P+Rx5vgD6MsL8ukV83DZIV3uaiELnpDVEt2EvVrexpkNYKY4A
ubLLGx8X8VJvoXdsmHIAMtct6clSE3eqB+jUHq8KI4BMGPRLy/JIbHfGnz0Xqv1bu8hBPea0Doow
jKBooALYxsYcHs8zWz89/IeCW4hau420LxB+zD0nYnIRX7mK9jy/xxM7nFN7Z02+A7SPMz2sMJ91
XbvK+A2HaOJirwWOiAW0cZUOQmp+KvvtnK7FU6Hh1yFl2fvJFRdgJnEXxVbMEzMaKyhoGU2XQF2O
H4T/ySWV1JZNJhMT+/OtNsenkFxFlUP30jg2vZRlcoyA1JcwECLzgnOMmeA0OCUWzE1Uk4FPNvsS
3tvfRhBNyjNIjejImTC7rB+FqCswSNmQuGpfmoIDosrm5+3ufQXQO8IxNVZ8PR+0UK9171QhcJcG
JaNZ4Dh+P+BknfAr3HV2B4UOxrsoPIXJjWdThXS19uzmd1aHgDFQl0KFiXkkB7RdnG33behJth2F
EYZKLcokFrwm9e/05FleKCKALfJPl9FqHnlyPVAbT6l981dBbWXB8hKXwXkotE8xPZqq0UUGk0En
E9h530qr5Puuexs3bAAxcFkwPLDq5TjfBsD3u2HEyybXbqZnQtQsrPIzAjtfWYsqHDvqh2HTgqOs
4mvYCLxdwLjEzeiGKubFs7386y3RVMziKbTmRa1yF/v6xqK/8+5hqPwGD9uFyrz9MXjy8xE4aOdz
UxZJSllCCs7EZy/Ve+ZR/a0GADg1l8qy7HR9bpIWddmfPIZPI1q5QO2AgjUaAMcCEhgRnDXu8oTM
fHyQ8+Y0nXhNVS1s9KsHx+NRshY/Ar+FJKDRiqI/ifW4kFSqMIEuX38qJqN0TRjT+dwiGIT/D5MU
d0SanVEhcYuq7Z40VaZgyqNgzz9X3rCzPI427UDrigctG5BhsEhXA0QPfwJT15b8hwz0Qa7i2y0n
IpmydZGaTqJIp/aHAxTTGTrg89SwSkon0i6Od4YfrpzdzwlFA206E6yx2DaS0uLmT7pILxfvRcrS
wVnYhA4elcJHo6kQ0am7L2HPGwJHpHndb/ZdKvF/Yk14PT0Lm1WUbKv14GLOC8OQ9Ms9vTkogbKK
m20+sozvmFXLhKQpemKssuS2e8X1beqs+Ro2CWBmVglTgZGi8ti8lMXXxvvPrP9Vr3128MK3017m
Uim/M7egVUJ986hEp13+1v/Uw/rvabzApeCcEnBWGp30TsTWq0gGwJYh86n/CNL0KgvLG7Fv3IJO
bqHFE7//1iNm/LTNzfvfqz+Y4L2EVgG/xtYRsYj3MhCO10f7eRTSFF4Ik3s0FaRVkEUK/Dinbi/G
XVvfEf7WQyLLj2se8wacOOeE2LzuvpFQdZddLN0drjzGA4Hf6kgp49DkSpRFbx1yu+Mu7jeyA3nV
CsxIadqsx50yF77IVgFlAjaFlBAiADpvOQrSWqHgIV5azXSfrbSUSDGr/fJ9ygT3CIXuFJjU4yLW
UgCOXHmfJoGp7kScnhQrbp5l+EIUIi3bFGf+S1vuHU88wyBHhNlSINv9XiZp02khIHl/9pqEA1dK
608/EchbHnuh7Wto9lcMiNZU3+BzzXXhc0AB73k0mKGuSo/Gr9Lhx+JqOxNbFsELRYAJZFqvUd2Q
sblL8pXrq6QIU9oeWQ7OeES/OYGbX3kdpr9R9Rin0r4fw2prywXrvRnRlnJgk9a0zfYVZYvtbro/
UosDx/+iPtYv2Z4q9QPbiWJe8pRb+/wO0G++IEZtTFu2Ik3af6/iP6u+foo+h8d/Wv38iVm/qtHi
3npDwG0eDKcI1Gi0sOCNt2rsiTkUaBEnbxAMZQ50WT7Dni1wph2JNAqujZe4OEwWXz2mIj5dTaeo
FFKNf4FK50DbbTy3tKSWlXiRji5IEi7Bv5ap6r+vw48xINkUWsaOLkO4ShDB7M8ZrQe1OJKTl9Ea
QOjPJ+HwQvkJnRo4GaLh1lc4oPiR9ZxGiVhK3UYZ+bjqUSioiNMJSVqtxJA9tzuiQad2uwKr4s8x
UgdCxjyhkh2854Fwa+GfyH3DAMU/UQfS4yv8YPWh2OvT7g/VB/WqJQer2ESzmaVzxCPQUFD+JxTE
X+JYoZfN1MsSSNTCJbKCqb/tNPXMEcPmrupEbFVqYMU3EsKF7HDqdgXew7hHIjDZ5MbDRp9kKj5D
oh3gUU+iO2aAoI3u1Z3/GzzQvdpgAsUfCoNjUGddgPQxfJsmQTDarelglqzMTYA6y4i2Znz5sB8M
9xysEmuwZTLRRCHXpKsFfLGuxIrRw+3ZtMN094IhNu8cSBtAzGP2Nb4RcWRMLmXU8tnKhIOtAOAJ
e0vlDe6PhrbULGQq0YifykKWOXdGFH52SWdsTkszjb4d24KypGxtPk+8L4ehO+mnQaKpXFeb4rt7
lTm/Wj/xt3J1jqcCj+mdN4kR20wfj0Ji4pTX6WDLaPVLFAO3jbM4CJaAHkAB4XtXPi2M1U9psA3T
IaumYr6R8oXw7/3vKcIzhDi95SwoeLopsbldBDJpOdypLkDr9rKLikluCtvdf1bEvbrepMSfv1CI
H2nyDA2f77PTV/URLkjwVdAHmqgN/aWqsRk6jH9lM2SJ6r0pIJZi2Lvq4FDhz8e/SUoEGWwRdeP6
rOKzr2Lv6pPEnx8yueXE6U2UgNwO0+jtxfjU7tdQnAA8XbG1i5tURIlU3GBcvjYwsrTTXje8qxtv
qf7QHRsPvS+WNBBcHhnEr3coFKWz3p0meUNmyP+FzXIs5ooO6UIlR8dySOXDwk/OcAVF0PeKu/Vq
qwPmkOJbfmb02VUlrspemZFHCkiHl3QIufN40U6Wfp5eKJ8gQBswpBteIXV/rF4rLLvTd2DfhV+W
4h6+a3J0Kxmvt3eEeSguYSaJiiD+52bkOqYZXX0R3UDv0EethyhWGKSZ0goOnDhIz76Es15aC/bH
wneylgvAlgbn7R+DUyk0pQ+I1q5KG6l8OnmyIYfBqtry0IYP7G+QOQBJlj2rUklxQvI03rku0Ttv
DTYCLw30by7LpaR5nZMo/14CrOZVBC77MCT4lznvDGUTKWGinT+BWq33HCmjVdC+risiraWeZWAz
Woc0P/myan6LlukB/Bi88kO7EvHGcr+xU8uikjcl799Qlzqy2JIGW8mK6d+bj3Xz/c0Ql1Cd0JFo
ouEOhSGbCBgpDtY87VHw9oh75D/ye7ArMhS1FI6EV+2I5j5EIvG3z22dfSwjiU0Y+kr/lAZiFF63
d/QU6x7xd2hGhvhGOfsHjzIILJu0Mjf87fVWPYnIPEdHVgOMMqbT6huvAFxhuS3qucQPef4BmfZF
1kRSKopD9b5KNqLXGaeguo2EyY2hur6AsVidFA24lOXtfzO3LiUu1EukbYWaRcZUSMJeJad/VRAg
cAVNnfK9f5hYCsGk3uugKt0e1+2PuCc0NLB5TPEDir/BLXv3ubxpyYsvLUexgWOeGZZHjLI8Wjpc
LjpzFXmD3WSwMUYKb+SO3vmgwClg0p0Yvc6UWghxqcBqnbjLxIigONg/CZfNS0ylpWlzSC5DZq1t
b3tcBaF1IfbB/I66g5fU9mNd8c/nVbxOKKGfbrzbwAA0inZh7b/gAEV5p5OgM8tylK5MqboCvs0g
j8//xQ5iF3tmUMtc0UCVg0eyS0HYF/KZ3kI8NBlJ0cWel7wws2MtoCVU44hvx5xJD6mdWGuzeb7x
vtj7Yx/KNXLsndex5EzUeyHlt/XhaiiT1Fy/vQjdI/U1icMP6GijdFUvHj3axrXy8ktQq/PIuBzH
O0NGVQ3bw0ETKsdmon8Fr/TmwUGtFx2EAptsZredZ9ECh6s96uUPcFVgk5f7nIddoVg/H8F/xFQu
0x8OGH98Jqd6Bmus80uqVsQUQDm1gYyzhao4HDkdQZ9SkJ20cit30ujFv8xMJKrIAcpX26VsBNrJ
NuPz9vNcPK7bNo55HPMRcDC/Cs7Wg1CNQ9+g4+J0sG0dEg9aeAroPFZ6mIE6eMag67EtSYpBunfn
BQZTd9WmJ55138ugStzQ9E3Id1zbFVAQaSCgism4yGpp+W6Db6hxa4W2yzj3efPF9lSlYT1tJdZZ
JRHPNk0tJjCBvqzWKlrGr/uPrCacFMUmfn2lnS0SD0NIndfq607nMcvJP2tCXSu3cMo61Y10OFvH
zMLt2OgiF74HOyX7JcKh0g1WhKzkMXl8u/uZhc1BKasFv8wDP8KWbWhspKcdeUkaFfxO/wAW/Jha
4xcO9YNbL+CHQplctoE5q6qrbLrAOoFKQV5J5iYJ52++sjru8eiK3X0yC7NRFAcpQ/0VCC1YOhl2
0ccLxQZ6lSTherzzXAC86myjR3Ju6SzsIcvOexhxhV82ma/FOsje27ydVpFzcOC8e39vyCGuzJR6
BiD/blyebSIi2FVhNWNyxn2KavYqQ+sLBw+uvaDIsrXmTAqHnXlFtn+S/CvzIi52sUy0DfqGE7RY
aH0B1bZ0TS0esZItD/QqopXnrvUU9UMmbCJq6sUyDLElK+MsV840nJDx15GlrNPPVjBw319Aoa0F
qL+dgf8hLvEO9lg5K+GcmFD29gmbjx5lqE5IZ88pY6yR0VugNlwBTiVSIIuZmKi2jLwnWRJ0cXW5
/OE3s24xOfT++o+tYhC/F2raKBmjtItclCf73mecDrq1BQpRAzBn5U8WzlkxLvLnxRde2dAoCFg3
oVF3sf70ghqhaFSF4wvlO7xjwwfi0pvCXnMFqHO3uNXFzy8Vzfky41sPZMkwjdwEX2PtqXubY70Q
XrtVisLq+6qcvbMC5Lq0B5aWHqdqWDlAj2BcMsvVoVQMr1DBnyE4dpNSkYGVgrz3mXgMIUYaSFk5
oJ/UxvlXyB8a2pNnM9WhMJy1+Q36N8T+qZ2E1d3PEfMYVm+0wPznid4L98cF++hRXPSLmemiFyjF
2sx6o01nBbgstBtuxZLF8Tk6mVLMLefDRnY/ghLwVvz0JnVVkGHI2cTHjuwjhi3+TSrYZQlqGxIG
vb284YRhNaMU+hxAMPPcrvDFfxHi/8InUN95lwlO6Q6zCtr/fsqLmt7NTgirNQo4RQNZjExEd0fN
o/X/QVIFHd3irEQRsHClNKLrt/5vLVgYumbWajbPgtvqJDfNtPxJswMC1gKxhiE6EpntCAqL4yFr
/fGV4JoTWUIwb60GMxmGmRsnI796ROdbSUFUYJZxfKrA5uJkH1p8OAqCFdhHqCcJPvuogXj0Xzha
/XeTwf/0ycRD1vioWwu33ZJZUG3kJB/g8kHMUMzaXriSNom4Wfx2MtlIZHxl0mtxSDecfnRR4CvD
kC4ChM6yWcszfR05frGk6o1aaVxCJUznhMMcBX6Q8eKFIbXDkTm/G6n+a/Oydz8icwxQODTqp4Zm
2Vq1ZQO/+afjUQOjzEJ6kTJCt91RR3KMgwlS1/ZV6WN09eN3p4TDqZn77nSGyxj09+OuUhYtl4XZ
lirrZvdORHE5Fewr4XVO5tcJCtuFerYWprGpuqdeYDrlkEyayQG1ooPSp2+W7w06WnsN2mOzxDb8
0p6hF/eNumBz/qv3+6zMWbEGYFls6xgvwgMRcV+EXjEHeCqOP7VjV4NVLBGnV6wsleMpy93uXpQN
PrygbUDj1dS5JvEO+scC5QuZbKCJ9Yz0uFnbyPelyLDk/KxhJ7EFOqgPLXysa+Mc8S88oYxv4oqg
NxdiAs+G0UD8k8eRGhSJAkxQya3AhSi6ViiT8mMClapUxnPFd2Id/vCAUQyozqVc8H5iE4JqI8J7
wdnZSXGl2r09HEQDKUzmqL8CRA/83pO6jukASRK3BTovynOK8wzIvFvjVGksSDVwlOLu2wA61Prr
XATsfKnoYv5458+yw1mQ+0s+y9pGQeReyRlju74ND5RQLkhcj3tG90XjcylHSu/JcxpzdwkwNvef
ceivafBDASMZr3Rt5ntbFTu8ltxf5JPPLoZgd3scAxrYTqF3512guYStR0EFedjooi6HCqSWg+AO
2TpTuIsrckD5lDmjA3ICWkXCLXJ1/U03ppGttuYqyZzAjqF8gEsZp2T0ekxaLTEAhvforTmzTnBc
9fZAPNmodiFhquo7PZ4/4zqX0qpS4u+3KMSeRvbLGFD4dZi0i0XfP5z6YCYovyp6R8twyZioEnJs
kO53vts4iGYWWqCl0+i5c2CqaAk7wYLyJ6ny3jAPD7rEg61ln0s4lHOalUjp4XFLtNWtyS5oyLm8
vzwvfYo+EDajy1ivoxqouvV4cWmTxm/Bb+WcFNb/MKwAcuR7sidZEpyLg2h0kd5qUeZayvels4ET
MluLWx4+CuFKbaKRHUgK863CCroNxJWSVlTYxTHusYU09JAfB62jhyHI9WnXJ4J/g+0kKb/Grh/Y
7EML266gNKYBsLS99fLFtGbpFqDM/hf+za9XLFdyiQ9pIV4VO/j2duC1mUqWnD+ihWDwG8Aj8gvJ
snc6XhiUHvF58CFBWxM67XoO+Tmp5zKKBiMgze/UBDhgsZvQs+1Lc1rTWsUOkfjpOXjCfzVjMvCj
LFunPxDI9uRhLdY2DtRclp7cabhRhDEkHwqdBg9KngLk2c5BWkbHUXfKG1wU4mMnFWY42TP6x49l
UW9stCBJCsQJ6R0peL9Y08r53LE5J0R1inTZCDSoaUfnJDsMtNu16EUS2mCwNAgrg53ZX7tuM0Ni
10Y+pyAuDXX41onXOZ6kOLDeL6Kse9rN/hPXztJ7CyoV9vyPoAFbjfx3Q30ei3D9uOMxfpsQO6sI
NC3ODjN8oBcSoOA1z7x3WKTo+zG9d5qSfKBB8qetLelcu/dZ8e9fLdPa3EE4DqyCjUXlOLSOO1QB
ViB+UqwcUonFAUrtFtXYQUg8nOhdLfii5+AdkxYBh6oNo+a5ZyxkVp0Ruw3GLVqCwf362CrLCr8c
lMIlZfGnvjCW/YRBoN9Lerywq/2jrkd7PQmn6Jy1JPgvdxdgPf7sYX8sw4dlxXsVfZ6C8YLLx1mA
qnkmKJwLfpzmAbTZX0RN8iGrs9jBD+3+Twq9Kkj2lNclazeMSXElQ69CFokkAC9evZ7WfYCTKpyj
qyxgFb9rYEp4cYufx8+WFtTWxVCVA9LDKbgNQPYaN2pB1uueNIq+gmkBj6ODD4dLv/8M2Agwg6Uq
Kf3CYexr9+aHazMd0SuMYXL7D5uG8KByePUdXo7dg7fsMS2WD+QD7yvz+zc4kdYsg+Q+yA6AHGaR
uQkXEVUHKvQqDjmJZYeuGOGUWN92UoXRwvx8zqYsAjH3KHPHI5ZqiyyQZifA52nbhH6qOsBiyGaD
UYsmXwzMarfyzLLIv8imoz8u6QCd6mA2s0a7N0SxvZ3C9+FKaGNb3U7/4rXR4l9sadqAoNTdoybh
xFzX8phnHpouzRPfQOWUU38GtUB7owz+eJuaSyw2YIAX7u7IPLUicCWFK0Kf/FrRd/iD0ZTQWieW
xh9PPlT3Q+SYNOK++hlwLySZd/ZnngoqZJES5sBnWWnFcvNG8OAGKLbTZtkxgYzrEnjWbgNyx4F/
1Kg2I2QuF8VjbzFMXqhZILwdl2c9kIGZNrujDMqI87fmqKc+CWq1a1a4ZJT3B1hwd+CcODbcMnMS
R5xqaNrsAipApdcafIXNny/Ja1CBxNYsQfKwW6PPzGOYsWCbOdigT3qjJAA7mjxrqVkuIvvOxc4H
JlWntZyMvMgpF0+1xNcmdqcnOVyzkUrPVCnlTEUJKXVFRN0om1MAM7gLv5wpARxN90MzAmlUCyvr
q+hTknS8qM2c2LJ05vUSDOenUuV6Sfc4F0INDMKWOhA5/8+qY6nAAguWW23ChktZ2Ov1DCSmN4wY
5UpOyyQAT9MIuP62R+z/iZUai4ww/gpEvFgtPRnRyTkXltaXMeWrl8eIiv3++4OptAV5V0y5+nGT
WbfGYgA8weRqgvFIf4rKaSVt59v6H0HpYGyFYIgPfljYTDXYwEfSujKaRrVRzswaTxgzyOWqyYGj
lSsfjgFdPbsK4kyX0YIogLVX5yOGqjDNc+Tv/ZnmTu4WTjbUNQtKyarEbsinOKIwAg44lU8E0wNs
c8nDmNkVgOWmXmqjgUk/4mjPcy4wnIiEj8+nvFg7BXPKWLR3GfUfz4zlOemSXqsBkfeGNOE1ECfs
RDhWJwQTXvmSHQQGCOr+Huw7KBYltMT6/3O7WSTm9E6foBxVz2mXlRd0z/wRsuJgWtwQLiSPE4G+
1EmNj8FCAwr6GWOmXNyJvFP+XLMoLwFAzHpLJ6tZMpDVLbn2/hV6spg/+b1BnVEVd1FAS4Q2CEDe
IFIRqwHIvIVLuTXOltx2cciETObcPI17H8CpCVUSsLiKIIOZJvGNh/E2klAXJ3d6dXbWKjA4rptd
CPDz89bzr3MpjPfiwx1Wr7BP0LU/Lv83I4lszBnF7Y96Czjwb1ZEvTMM/FzRYD7qnmGfOKSdhRgt
VYIjBBoOMrpfquRNULMtcN4tfgKV0tR4PzUHMHU0/RFlRZi/VGK2mrTZ92ie1URbs2SSTFOxWrDq
hQGeky+0SciNC8Yxf2O9+AYGrA0oEVN8oz7e1/UZVlnhyO3YNHxh7AlCR2McQpedgrZM5kn6g7l0
KRMMXfjfw8M8PqcOOWurjOOx5BPPTPRPqtiislcnRrPkQYrx7dKH8VUoIir+Zq/uSDvAuBE4YC4I
iSNXT9xQQaoV5qnYTHtKMKBcFPO12OAIKO5tS68YvRh12hx1mByKDJqFJ4BmsEGjyAcJH6dw6cEb
Tf1zjEYlJgFg39ZKjt/PfBq+6AQcUvT1qMdPOkU2kA+5cjv78kQuXKmi8Yvx6xeMHv0S3rwAlNhM
3VtWzOjMeJ7qta5PL8doqyAwwEvX/9g6c4fP+M6+RALx0BFkxsfsdCSBSN31gdCH5RQ4UgRKOMju
XXmeANBAddXAWLpePeIbi00sHcnzeTmk6hehsQgjZX9oEbeGv1IQGWWbTrZ6l9ugyq88T2fJ9yCG
LFVbATiyJgU1KixH8ZzUEpNM94gdexwU7L07sguOqH+tfS4vmeWjvRWYbAeBpIWXhlvFwAtsWSwp
lCsv+zQgwNtykGkKEqkiTs3qxQ0RxCER6NLZpWKubV9eTxQeJiHR2GKLDfbdy1oeN/Um+KVl2Gb+
oSdlLC2mfLSYWm2Me1HEwl6Uv8Y7FmeYpxVXYcgaN3nkcKkgnfdJWwB+9L1SPJwq/ud9oB0G4NY2
k5sO5lS1vPD72SU9Ptf8/uqjjFy5ncJLPfduIHyS6wXwkbCWmOWG7XEaNScJWreEgYNvvyt8c/o0
6dYfmWbL70yE/kJd5KIzsC/lpOd3jEGn5Hffo5fM0qGnH9RnTmrDfnAl0rY1D4xpmhX35GxWtNHh
O/RNzCNn+iMXxZVwNAlgstErZgPJfmCcuIfwcgFZhV1qfhd7u+DS78T46IQtK5XlReH9RF5/oSMh
7IyqpWWFhw63w6RJtRv0DIN6W2hBIVJGTFmtBDSkidjRwhSxmAj16+GiP18vlNU9k+zjeW0aCFnN
sgR1dIO9+xeIMQPQ7T1t6JMW7E3gqtv5jpPSfiYbDwLMNdDNxLBLLM4Q3oRQBt508bQy9dEqCBW5
c7VcBM5byVvDY0C9hAXoxO2XF6LvVijrjIpAftAbpyLPQZXrTP5d0SlCCcnvloy4L1v5RLJwph2L
NrLKtsGcuILgZ0RUorsYUgk+uqmmgtDbPl1DTRpTuxAabZfe1sni0QWKOoQLn3LfQMhnKkiFjwKP
hRdDoEEJFp/B0SArWSQGAGs66d8MZoPY+feufW8rzcetVCtxqtoucuuuEGtXPcP7giOuKvsh8ZBm
JGAbFvzgYpMY08nbDMeh6El1TXkOA5om107qF3UL48pwg9hAKZ57+yQV47r9+MItD7f7UJcDdWd0
u4OdSZf6ror6P5TSyxOwoTOoU9i7T4dW9EjErDY9BSzgKg43Yu/gCO8KL9HPwUexfNmMw0gaTYO3
CfH+oDYpbxGVTGCbqMSWsjfaonh0XBsqWEQ2PsfRaq53O2wCRx5n1adxmRcgIvLdl4NhxUHvonMm
vrWHn4b60PxGEGvshiSWKhw6Xfe7Ynqd3lmYFnYYGrfnmjTGZV3QDOUDnblgf2pLgL1MZX4Dla/U
8dr0JDdhhbJ3aQD2HjtaOEUo8FAdkbJM/eCJrd9tlFF3urVbDWtuqjfyNqlfzqs3K4blo5JaumoN
QewYt5fs0thzXGg45YUjDuP4JU+Ym5yx4z/h0lxA4InpzBYPthbIoS7OyavdSSD/FFjKZuCnCQ2y
r/Lo1+8XoEmhSKBu1y2cO/I9lrBtXDJEEss6WHLAqCzdSOOf8AyMTRGhWY52JdrWvvXOl220d49n
Yf57HBLw2S+Ilu946aWztsRAzA7mC3pbgkezSQNBUURQu6WVNy4dFunIoRevmz4ITApziqBqDLu6
ouPTPgYUHuTnQ3BWHLAPyDEsfkzQrjJpsXHMmD2J0BJz6w2i3LBZeL82aUhSl8bOKeHWXVvOzR0U
RLT/gjLfEclAp1DO586cr3fGvb1jYRgH76o290+jthKfJxKwLgwRBO4rV7j39Ma66zUQHR2hsY+v
CcAdOC6fUGbocxaa7wwGJ0WcaAcpiEZd5qm6cT5UaiEJjRigavwbL97CIsmDUVYe8LUJRr4w3+42
Fvz3r6CaItdHSX/ydyNkVK4jWlCigabKMXA6EM+0NaLCYhiti3mReg40IA5G05zyYdaKs9ib07fJ
fSXm6K4ikO+S6WtacUAQuEQv5Vz3vmA/sibkvf7JzaOX1DAvACrE4MMU9bPUsgkQJMD/vXxaFbcc
2bificejb9NqM7BOa7/BfcaBj+pb41rsoIx2/llCJ0ydJ/KTKQWL96HVfmEVpfPDsRgT5HHpGZNQ
FQfL6y3ZzpYrgBa8wZ1I60KL38htOor9YO4N3N+fbWB7hC6M5uSBbVF2w7jCGNlcApFGzrpA1hRO
vVzNGBgj3u1K7ScuOaLh8YyonpZPsAheNgRjKByEz1qaXvpKnEJMi6AznxHwnCZntaMQyv1gOiz9
vKnn/vpAgVx6i2uZ1Q8TzT4/uUsdtpjdq3mkwyQC8yoERPE2n9mTeuvMyCB/3urfeQeWHRA29/nR
1vfo1rFkYcgBGpgVVThV+Gu2PzpnKfJFbmPcY2VB+hnpngsrifwESks0dHdbWJEZkxXP3NiiKywh
vLA/MLL0guXKx2kN0NgjpQ/VAlweYqTO/xmhu0yJtjqYFQQUzbMBj08dzn3awMuwumWQ/Cny6OjX
ebk97YsEEAYGx6yCSh43mOo0ZqRTBdY09+GzFaDzVcCNi+CdbB2MuoaPaTUlzTt1mQ/T+cSOFdVp
HfPSe3iOeFcv4r3X0AEJKu75gmbqzcjMd5kzmFp9eOmrd6x32c3xBELBNBE46Ynvk0Nmr7fhEQTt
rp5Nxg5bzFBEdbs/xL+DEnx4z3GsaxWyQkiSywerOATfROhRFdLjfkQdQZhZlw3EsQsjV79j/rtf
eb3p6OdLKSpKgPIrqc9YKZDREsn+SRoAYSAbMOP77xdkph4LYAuYAhnzordddBIgD4VtJnCO8lhI
nVkG6bC/5WslElt8c2uIH51SA6Qe0vmlKLvDIMqdBzxOvjKqmMbhf5rbsYzJNXix/TGDpsPGMIeW
HzHVLlrAl7iWIw/ZUWt6X7IRxJgU2WiatMbQCFO+1HFMa25FOykai3jENFDZ+zlbdxSezcGBm90M
q3U17niW9or8P2BxHCLLge+d5W2ACMGMAjNqyZS3VuztwVa9rZGNq8l8yBQUyoh31zqhaJ9QyN64
X6zgK9SAPiK+M/lu5qoyQpxpWEOsJODR1iIxAORu0p3Ap3ULKFcVVSDKZCNEaHyvdveLWB3qpc/s
sAQVQN72PH4bKEvAmFTsn1l4UMWf3nuAJ7Si3mxJfA991gT34aBFZSBJY5R/oVzXbWSprs3sQ6ST
NVyNkYSlmeVpRXtj/tAoCv8mknxukk2+3RvsvMCcu57IuSanBpDBo9zUsMkEIWZGWnPZjYPVe4/b
F+mlxfXhnmE46vEyWPbSI/qVmoN+9BRVmOwZpvIrvVqNSdu/Ocw4QpPY8qQYqryed/Yn/KxtJvAU
id1HhWC3JN1BH/5v2nTRxaccYdaaJRSIFxCszCG9TOGgl1N0CRzxT5bbs1psfnGSGoEePCMaCFkB
B5VeJTXscpQLAcL70g1V8zPteH69YWUmts8PW78ikkzBhUvvgcHKRmf8LuOBYPE9dYpARq78zCj8
ykKbsBPCh/mBWHDWoSXMMT5HHKNushuVQQmAKXLlbcYnTT6vfEIVe6CnJFKBzcFWYOXaWPCNTIIY
EzQml6hcYGo0UDOHdIxUYV2DXFach8buoF4AwA4NQ7N4GlzF2DTHxeTimvIcfWDscIsXzS98UakB
h/VcGVsYqNSKUc0o+jPqUFBqTljAiGwlMr3THgpU8Fs9zdwvs/YTFvGQHlZHvMbRikp9ylKdHr4K
/JppDl49QvyCaZ7IpMsffOW28Xeli2fPc56ECS2BycHEZACnewRmMagZEv9zf4gaO4VEcyE4KutS
+ozE/P4+oehRwKYwjuXTrwYzfDLlNqQsWKAzAgT99H/+lGHH8vK0w2Phd/4liI+mHTNG6b367aOl
eVXpsCvD333Jafa+L9r2e1INp7XyNDJjmZi54nVr2Gp+vQQBOHgD3DAMLrtf9xpemm91nY198YKA
FmpNbVe/M2RrcE7+iFTYjN49ONiZhWYDD9KsxsBTDOOdmucCDBv4Bj6opw4jr9DQZ5EKRuHzwchn
s8dKLqUIhV1C27cU21RV+hkCPDczmHXawvW43CRUMUWLO6XpkozXEziA/RMKZRkoSlw5eESLvyNa
zM6yYhgvtghKnZZHPqsxThFXH3H0h8BhlhLyA7lCJLF7ml5LEdoz6iROvmXjpwdXttmaEP1vHjco
7OxpekhwXhar9Nmzxd9iUsseh4nA27/30+HgNflrK60rLPDjLlkgPKzeqMFss4szcdCXHfUpnVEW
hnvI+7BQcmVSr1A2kGuf7M4PKhKysJqkmINxDGVoS3X5Pq3nngQrf2Db55wxoe+52jeGI+Uu9RZn
RHktUgeuqZ9yQrQjBiDWJ/OXOYqLPGarVizmv5jJ07YThJzB7WEZ8vd68vnXRt13hpn1GC8EBk2R
ubyQGZbXDsF711zbyM24XEJM2ftG5og2Mjit5a8CgaGAs/33K+wlssNE4vJAzBHb4Yq5s/NBhusl
zrj5vbLaHzyhjc0jxrgmYE63B4tUqyGoLtg9YWfiNeBVAa0FrvigzSfzZ+tn2bxjWAgx163EIKZc
Kp5zJtMrj3IS6otQLgek9HcfjYSbC7/GSilNg4Zb2bb5PLUOqx5dgkUpiGa1bj0AP+FEHOLhEtYt
Fl77rC/bwPM3XjSAyxdSLDnKKPpgQVx7d6VWv2y1gdzivn3qL3O9XaKWLRBDjb5OPkxOX1U7G4B+
uGslU8PjzP/ZlX9YlqLSMpH23lkvCk51NGKT2CrPU0wIqam7Qs/qDI3XjcW3yRuu5txS9dsAOTqF
Ys7Ff4r0AEYUFwlnm7HR72DBGKEcSOUMkkN1r6xwkFW/GyNuEQVYkvbzpsecGbfQj9++xcgx8E6K
Va2kFdn//Xsh1WVaWD+haKOWKXpmJwFI778GY84VVO2JO4H3oDxlqB0HEcKonBm5bUpw0RD6PImR
4DEDkFt0Ym0cqV7/h5DaIGn3D/qWOmWsy/8K4FNlNYeUfLniHRFRGa0AGVt42LLpbMsT18XNtbP9
7/d1wm2uj5n6NHP5FYG1eRycHmPWiZ7dP43YMy3ssH/g9EIx82R9DK4LXeNwCRyhyZIfYDtCxHAK
RiYbN552UZdB7QLDlCzLyppUFRR3L9lnDVvSboE85xcckVT9kkObTA3Xm0dJ0DRbz/lhZrce8Aet
AFWkShPAT1Zn+kWbwfdyYPCpUNmY47ynVGO+V4XW9wUB3LGYXZ1wIA7Dx2g0Cx0qCGM1zECk6zji
NiolQaq/FW/uGTQJvI5SxOHj9ggJxGke767/B89oqWN2ehyP1xCRAbKNu8mwHc7jeGZBWFKBUe1w
N2nmeVYP8AaI3PYnSbSFznAr3SiBoxjsfFu4YCkKh/Dk8MxEn3gzpffp7Xy+8Gkvb3yTOhLd0C9Z
4NosHmPBltGbfWztWhvnE2f4oJj76SdfHAD8olgEhVQZlkMkOgn6f9nHZZpuJ33bF7jYeIzASW2X
vwLWvKa6z8Rgqh/buGQI2LSVQue5SDrGrP4Yvxl+TTsKSQRazL/W9r1Ok/wLhPSEkM94haEOeCme
L36bqJHVPGpTebnT2Rr/oVKA3hgN6RJB3SoashT+zAhoaW1a1R5KZcJ7xOrT/DciDJ2ohNQVICJs
5ZdmwJLZRneSL/azJMqkNvU6H2vMK16XJW0x2BFWTS0+KI36dFy664OOcprQTA3XnyAye+49HLVE
asRMYB/7l4TvrdxAaCP97qqOT6+eQ7ssbo/utX0AoZe5lQIh/ODBZgdjp99vhBvMn3E5vkw4vuPR
VGS+dZ/Oajol0cAgN4GwZvzi3qSMMgfHyYddG+S2EyBXE2qyEeqNFn0kZrrfxRl0wTeRjrZaBrc+
nsKTm913i2vGHJepoeyDNW+/Tn8hB3reKQQMJL2BstbA/bJyjHGDqWOOTpbkNFuv61lzOeDFvSL5
5yTsr6rgC5Yf8ItxIFj5VcBybdWOnqlPFj/QT87xLV5LYeueknO4NfJMhgVDgq1MeeEim1zmXaUW
HZ6lxranZJVFrvrNstIYYiLREayGPNPVyu9IOahghvsaj/6OVPZp+VG9nfyoH9BBBqGordiOx9uq
e9PNWP62wYv270//kXEMilSxOjT88LRwpHDUFDHqnYE8ic+gk0Zrc6qo9PgAX+ynNz1FcvoJTX6S
K5BbSVoeE8L+6QBf4Yu4L93FL0AhQgoPTuRvwE9g8X1JPfVpzF3MzfgHCUM/qqA0sGsur+Cq9+2D
dvbJw2BTfWD8QOZLnswWlsOrWlddQOAOXtoEZZPKn29AIICkfCymyF8pboEyHfzmdBo9tt6Wex5q
G7ZzoPePZnDjiS1k9xyYCSa7vTUzYah9xaUJjgkQ8DLih28FbXDc77V8ELHx5uxzTmXORO52rDWm
TJPSdjD6hyhErY2+adyXjdZuVgpw/2LatpZSLyqhRIxovkpWiVfgEj7Eo39kkCKEQMzbR+6mvibd
behp7A/nZeXIIFukN6V+d7cLVG8DBKVryEOMoc1yTg9LEe0DSHBMLuaAxYa7RIiHgAq9a5YAvuyX
2SxRlkpWn4sIvIUv6sAoOe9vp5XQaqbxvhefvxvSOm1qfKfYgbpxJ9yeZfPWH98NYIQQXZMzRNyp
c4+tKE4MGEisfjwXb7N6diR43fiD7f5akGqhBaKbS9eNTLjRbUzLMwQvoNBOr0fhK4vAnvS0R0wr
kckPcDzGdzVdCv9CBQnPfo5Dy+2IxEQ2QgaB7R6cwe8VChlrZtI0S/aUKzOr3rYtTKpgADBZbI/Z
JGfZ7OCZwGA619+d1WCrAQDAEVKAum3cQ3Wag42reIiFSTDttcW+ukKcgd/s9UNbY2c9J2wDipQ8
88M+GIcEAGtKzawLF56d1JieyPT0FZFHS7PbYLxU5ET/9augDgHhkSw2uf1DFtCcBU2MiwhuOz+Z
D7iQZmut8RPgTeiDvZkuRDfWWgXmmntOfzt9gHqH8OnPQ2HZpjleNRmiP1CLHTqnQyCYQuykgpb+
HEmK4V0ILBKJ1MOaUV9P42j6JW6Q2yMvu3KRcghrE2+7ybWWc+RETeMquIxkGhYup0RyzPKap0xl
bVpXD3rfXZCGvGfYMCqpkvKECIQiVEZuijYEzFqgNtd+bAATuzdP4YkmrSTL3i46WsRbUY+RAToJ
gRrjYYObnixr6iGx6Q6YloDF11PQtj2toyaTbB7EEBfzdqaXAZnWqvHLEYUWJPT7gPJxfEe+35V1
kkq/Jzwvkzpo1Ger3KETj+J+d9XdyMkBkcxWQLadRRRzSnUN5mfFwVa4faUaEilhiSTeYD5ZAJME
OouCrorK5laoQZjD2yWapfd0kxcQvfYp220xmKrbteWY5HZpiB7qr+Vo4i1I5XupdJeH19LH4/Mt
TrkYr/1khdVQkvK/FkSF7RapoSgIx42NsjmluKWAzLrpEU2+zGw/6PNHXtgQaq9IEUEhEzd3dtyM
Js6eB5i0K8uMpsa6AXUDfs+HR+PrXO7gTecSYL7KgWMccFu7tpF+nFyAf27kn9w7o3KlSA+BwCtN
kTH8hdYSLsDFQIlErslezGgbJCD9QeLhT6pqoRoRvZQxo8RBpBysVpRjNzEopN6HBCZfL0lOSVd3
E6blNOS6c5rO0FUNdacSIbjrYKpcLTS81+ITRI52i1I2yq1HsrCDJOkxvv48wXQz0P38TP8VXhHS
GU7UVVFTW3yTt4iXGJ/MrczQtUTWfwiQAnGs56VPZ8CwCbu94820ArJ4duVdtc13W6Rm49tSkCZE
fSbpIgp85ld2cwh49Gl4N8dzCMSLolFIJ/G+GqA1Y1/LVnkiWhNSPl58MaW7TR7zOYagTl4vS3+B
q7v1tb6oFvDxCd4P+OUkMZlTamjGMbnGB/TfPnRGK1LP2mcs1vmJSimYqOt8gcybt/KyJDo14lSQ
5ENRH/ZhuVSH/OHEKH3cDzRPFrTkNAkICEHwVMfpZteOEsisfTWOsYlZ5wBZnxXomuI3MJsn/iqH
+gNBXzE6WcZdxYRviFNA1S6qwPZUn6Lkuf0JnTqh3wqA7xMZrjXiT5LcNvfyDO72LqbOfqDBLgiS
C8WYKf97fE7L44HzTR6oHfsqPcZ4WYSqs8G+iZ6JOdBab6/i7cS/bV2KF75do5qQXvIkrwP9nvVk
nqwQ5M7S2NjGQE0L3Y+wpbjMgX+u2iHinSp3wYDuA8S3yjLVW4atW+okE6taKn+C2CoCwet+ilGp
HD8UZHGH3mDZHanEo9pQPiIrrV4BMGW0ZlfVPV2v2Aoog7r9j0wIwNHsqM+ObmSYlPT3kNCQzj4m
Ue+BG42S7MC++96oXxglC5Twq/43uVS9dXTKWjK35GQDYJXl1aA3ub/3Br87eUTyIU1a22QCS0Mm
VIzqpa6gJw9/ejGpP5oDaDD2YiEBA9epfd8cG1f8w21AxAkQvwSfuPKkZEWMhIV6AHeZ0gdjqbM9
1FLYzPgnlV/Hc8YHnnK/yAbc5Vhi6feXokegDQeufOheH0AwAl3W1+mzTezk4ia8RjzOVUysnIRi
EaPedG6i8gaAbH5zMXJlCXDibuodeTfBrulYlPBAlE66lNCTFsc4rbow5qzEBk486TQzBBUnJN56
wEh1ulXstMWDlSt3QhP87u7Mv4weG8RiCFxvKv/ZFzkWfcaKad7W0rq6Cz0iGGnorMbMb1daq2ms
LO2aE48aC+w/eUqcxUTpFpHn99Aky7hwIBlSCBnOHA4lTXgSqad3XGTKH8/OUO1i+POgv83XXhkm
bqXWTsNnXVpPVRo+D+LWxd5LRQfAT1sgMQ/qp0ttaBgcQVsE83C/tBgqstY4fja85o4CXWKWvKWi
Q3gD88wFZZVHn+MPb0MImRL7vndUwXR/RIMWuGipPSAJqtPQwHBo6ziTdVF2B6ntHGgUxX3DcnMt
ftBx74d3b2KzQrfwCG8ifRVIw6+c4n2BjrTahofYKc0kA52fYm3oTcebHgXPyHwljT8okG1+AcFD
GiklcX65R3xYDdGBkc0I2R4YEmnm2aI8pNPPAMTufxzKkhOSyjQ+bViIJ7tnQ4Nq3gdvJU570aCf
aDBUwf+MhVL/NzmUvUn418kMm4mBQgJPA4vFn8Xu6wUDfSkvy5BHr7zqk8YVbi8orO6v4iG92f3b
OE/oacUjerfIi9Ex4iShxJeJlEXuU9CTnrHfDOoQUpHFhl8vKGbiJtOb4d5LyDwD8UzBQzajOEqf
6eQimKK+xtMhJcVUbnbSBYJ8VGZ/k6gO5N2dKi5xhtEoFaWw6YEOJs73ehfSWEm9LEBZ3pwj0fWp
OueP4ZSYcEzrinKkz63r3GzNCMaAeDpl9eFMG8byTgVO4yFZsTS4FgwTaWyYnY2P10g9vjDHWXiU
/YY+lO+D4xIf3onPgmxHyicah4cMfQ6vAqZg9OUOyhbwIfGIVRH95SEFX1ucYNdYJRJvrl4Me2iy
82kbpUILmFdc21dvu/0Zc++Pj1OBvhcnKGuaFkjBLPDXsAh9bP6fUjztQXtQp7obc0BgfnWmjdps
jljbTxnmSgKl0FStZqEXb4KeR2ajlTyhQ0vaXaPJuYZiikHJCdUGgLj9lMTkRmmGyGVwwQ/ey/kN
yIliZGwRGQFtqdkmhSMvX+2/zxDFJDUPlxh0QRdfTPM0iZXDp+PlpPCgd3dpCinzejhbIdj77xJG
hOmtj4qulDHJIkhHtMQCCKfLMiK1+mD8m1mOiW+xoeVY4IXbMn+luStOH8VfBV5p4B8SyczxX34u
OXwFE9bjlz2ZXWa7ewZOitk/tQ6s7dv+StJzr99l8BXR2RXB8NHWBGNQ0b7nvxnk79cGu02lJPp0
vkwQk1WzxBp4VjP0t3WR8G0BGNwT3aDv2Y6Cdq1KAYrLSBc0gHumPltMmC3poZt0EeK2t428GzTQ
pZG585NKc4hdNMtvqdZHsN5clmKIKdyuap5KuR4+2ZxqyyOV2/sesQbg816/WqoAJ8g5ItqN0ZsW
6x+sTT1pcrdk+u64ZTEdHW+VPgV4W/0sWyz86diBIyZJiCZoC6lFyTKoYZX5ccvX6LQdLF9zBlwz
7hoBrNKPHjNDbz8yfVnZ/SjdpQ1DtCCliO1YjkoDJHLtXDUCMjBACnxN21FRRKn5353SvMOWbxeh
8Q+4T1TdtGnK4GjZhqs8VLDqPSmzFEAdHjotGDeOgpR1HFcevXaGdm0A5bCAmuNoCOcUn8/yuKVa
JRsUkl/Ssljv6ofJvncBOtgVcec2GpMRvr+5Y0nXVoaorcTFGYndwuQFqa7zb4+mdbUQ9Y7zSW1F
zsdRnpf5QLHJD7vYC3UxZk9/xLDMy9EQ9sbqrZDWTatxso0rGXU1TO47uOpWnYyoUdykeWV16HkN
egimVc8Klsk4aq1wKDG0/lJc9ZjLs5nGvzM609KDNuRJmf9U5trV5+Yu6B+EScWt2GpICXe8XK4G
q/tajRyZBorh2OZX8X9dSZW8Ux28cX5mOmjPUsV+DFbs/SN/Ku2LzM3DM28ZP0AqumCSFEgDJHuA
DroA/VLA+wHoHggj6dKsZOf6YYBvR+8BvytjhDSzez//vkCIlAoys4aXTmqH9vGKN1uXy1hkXNq2
XX//j2ObDL5/tYwZcA9PXwPIFO4JtMp1LFpiwTe/Yn007m6bmFqgZhsYR26Wfcg+g6CVwGqWDCwB
yI9WXi11AXWhqFwwbm4E/CI2qwqVJtMf1JEm3dLouA06cu9rlA8u/vtiNxVNsWeAX7lqlIz6QeIw
QL+b/BT1bjZmdB2IBLok6UIOKB4Cn+nlbDKYaVtjzwqb/CdhoLAWLmDuxaCTX2tcsTcesf7Zi560
VR6EiRGNV2166CU58c00/kwMlLqeiQM5GALURnya4WTe4EXUl9HMsdA3pn/eDJWQMYVy+5oCKI0t
AovJ+vp++zYwhqBRnTR9ahrgxGUD18U6mOOj2n97flsJiVmNF5aTVkgPjEwkKMtJBb/9aVYeGQtl
pssjBWv6SFbG5r/w5yJjhx5WeQBzkYCkH+xAhZSb67oG2f43qHj1eZOobBh6XlVYIinXraawqBzo
VsOYflh11U1uo5XmW/cUJiyedZ/fMp3S8R7g8ZzZtYcG7qmLiJTLeUtgTT3JovTWtIO3fI9a5F5u
6GC+3ZU/iZZVUyn6tfSdb1f4fpXbTAaeZyNl+QHDM7og+txn2R5TW4WcDQj4JBFRPMyhS3DClB2/
Jqi2jUMcOBKI6u7ODLBqby1XTZ1ve29g6Q36ll2Vl1o0KgbTnlI1x6YmPxk/GvaYiOeRsdN9m3IC
+DjTa0JnTeZDkMwyROWc+hNmgUKiahPfYvr/2SLfhC5GYSOIHaAuj0rrzcHdHo5kPYFgiqx8WN57
qIDuy/2muN0tMC2r0ShWqi6PHm+3TXp0Tj0gZmAGoWVITfQ3TM1J4RtJsX7B6NxKziZKhKWqFNIn
TgLlOQI85ywTNEZHk4uwwRU4knsmD6Uey5zXFIHj4cnlHtxphkt35Q6hw52ih20ejoZmar+qvzw4
X+ptXGJ2y+s4f892HegG3d2P9Yu6p7TB6RkYynIcJ3a9c5ab8cccd9nvuOfW9hdSqaKMhmiSQEb6
dX/2GzO1659FGbHIH2yXrkNjUKTjGTYWy2i7iinvMBl64OOGjsnP5riOoIuv5H33Siagrwp4tOKR
w9qcHtt4X25zgcpOBNtc+eo/6V8W+hZ/dGp9F8LB3vobONJJ3MAiLPfpLkIeJ8m4tCZaIEFnXwjC
q+mt+X6XM/TmMPXaTSYdgHyhVHgNbWFgHFSXc4t/PH8z2oJOibXbh2XTrQMH8ZIS+GjRzbXLPzNd
/rimaJMf/ZosWQ9uee8YaWQkjJukjKmKRGVxvqBB+WxVaqieNGx+a30T+RHNZ/u+AX4SBKA1iZ2S
r7IjqoO/BPmep3yCNH/1M+Lag5qHWTsN02PaesJoNLpr2UPu+OPHHnokVHuwOeRODUgivmYBXn32
jdehyxRMVLpjooWJ5Pfj8FhMMK7JGv3ZQbsr4u07biNDJOTF5quHr4AdOQ8/QHsTqOV+hszJa8EQ
qjda4LESWfudEStSFKYJKdduTgvaYurnNsih7NOMccH7XAl0RszonBY02gzbgsMeSw7YvrY6m/sz
O9vsdWYcZUP2mzg/aq75Ph182A/HyTXC5ixSrigqiODLnbp2DCDEPCQI7pAshrtTz012+vhs89Ga
p/e5UUaPzp7vwppHgbSVBP94swGKbb/o+a2JX/WYWYLJFgkD8u3XsioVajx+m1mbF4Xf3uw4LbWy
AB5LVegnta5pOI/uKb80eTR1H2oH19Qi3h2yd8a3yZIXVPjP9JGAySO0it9FEwbOipQIJOCR1Ugs
03ziyoYJ/s+UMvlvvjhZ1beFkdPOMLZcqCdGgniZWBZmIuMobEv1TkUtTg5VZVwwJrAhSzDVo7sX
zoVNzw9r1Dt3nQL7ikBTVdz8JFmp/zcvEB7c+Yt7l2BlAc1kkdNXO1LrfFxaE3WK29lcMuP9PEpi
F3QNAnajyC2OxbtiPXIoG6jgEzZJuXX9IoZrgw7ydfRKjDKpEsVEyi5ZGzS3fGOrjUjV/QMnpYYw
DvQ79rDgqn9PA7xkAE3TF5nUxbSHdlcCqAy55A9Htxb7TE4usueYiZ73WaFhtDEoOi5JhgwCElAV
BUQtxq+UJtqY0cix7yy4hBBpg6dubjYk+tGN9rynYOLOV0LGn+0YsWo6YfoWQii/RfnVyod5wIH3
8OPsX22FjOi107Bde9K8LAiq+J+NpZTqysYZDHxH8948WzS/2U94SpXo2D+aItzN23IZpGrVMHAA
k4T7rnktfm9h7hHobYKVODRGgFp+wBO5x6szk2ITJHcNNGnz27Tdo0pY/VCPhsM8ys38P6nOxK6e
2whI2PUtuPZU08qNpUztzJIQLujIrw6zDsbcrEbXLhx03Rnb3atNBgwQqAJ6hSn18JjY79Usl8B8
gI4oEvvzD2EYA/1diC8ivp4fxSySJ4MnnD7Xa83Y7gmU1m6Hny9BsLJU4REgkaIMzdrpSHEa3OQJ
O+CAqic9qv5Mb5t06DyFPkefpYNaf2+QiJvltauqkJFLlFtcOzf4M20qu5OchzSWmHWsfBuG7EJ0
UxfqfmMlB3U2/Dx6IQpP/W9CZrsRXA0pWZZyOqtsF8GFoboej7kCvZ49IBoFu53y5AR2NGOQNG3U
ChhHCbWemnuOozBWfhJqyk5+4m2eRSz2wMCo7QvVL2Ns7W4NXDDxknKHLrQ966utIr+p0CzhRKfa
YxNx1VpHWy7mTvMFQqwiPxUmBa56nRKUPBsfttXxJNeSvSbs61W32yNuiPf085GcVFOwK4tukUk7
eq/SinwUNIJgXbxFzazKYH4eS4zQpjyS0dZlZQxI+sOII8L5UNzLP1hHre+NdlUfIZGoM0x/h7c0
Ibw5unCn7Io+ftcGpK6H6X2svFaBlkOMrCmz6nfwsL16b8v1eKDlx/xG8kM2GsVYMbWDW0p2grgc
Ngsi8kkkgdWn8u4gK7ysyNOZ6oOCX/RoL8/bpgXFfJX5F00QQeVlf+YEGKqygZoP44pLhRagU016
2RC4yjF8K1pF0OhCBKzRscWQu+N+B11J+xqRMCfQjfBoqfPnpXVxNwJgeLasxAHUZxKpvOAe1rdR
9YV1pRUA5ekvY2bdUKH2Kfswvm1SWAF7rZIiq76dGYv5APXFeVSJCdx4sWqKTqy9iCjc/SyMKESD
TNLiwohBXeQU8KoUqIeSdxll1+eL/5BbV1bt2jq7bYflWMJA1feu/1ItZkv9RYT77+no12lSERZx
JCX8NTb815yDFfSlUsY4NqXPy144J1fhN6SwEM1wkkdYu3GXkx1/jbSJ+dD8xBuaaC2xVcqCkxGk
fcd6mDLzEZ5DNAgv8R01NnGBKXlI9ffojLPE8w/cG0oysz7MTzbumIeIoEK7iOFFfY3TOdUf8X+b
ke5+STW6+uf8NjUAQJiAk2riEDMc3KIGUxXKGxEWZFhkERC2OIF6RqOjIisiKsXq2crqbJSwF6Qq
pbFKGDEt5Qvst9JbJrwQ/OEeFI/h+2UeFLF7ujHiw1ovc02cuNsHhGbsJJT9rdEvjw66sDqCagCd
9lsrddoC33dEzx7oztYw1L+j1C+C2dSKQZBri18KFSby/ZIAWGXbGEY2MuWqE60wUjI3PdY17l75
PeawBaveZTlFxRhnqcXxWdMyMJ5LTN5xyAYyC6YBeQk3LSN5+1QpT08d3qo7QplWok/3F8825KjJ
n5MCX98PnzJbmqgykxqObHurLlgy8GV0y0OQVHCSgG40hSp4r6CGnXfto6Bs1Z/i4acAr5E5Ajvj
SUUhC+VheF34e3T+JzE37mMPUn3w4Q0jKouXeweECHajBM+ERxXcr3nyNyb5JJl5AMzsuKqhIFKU
vlHnG6a6u+pi/vtjnyO8cmYOgu/iblPGTeGZmEXEYViT1+AFqiQ6FEXZ3BRYaSQszcpVKekezhS8
Q2Srs/qRNFGjY2WA2gWSUITEHa7+QWo92Xlg/cZOpnKAIX5S0waAwYuUAio2TH4FuRkUtzoOMoIp
osW5CclqoEXlfePhKbWcP17H505VKd3QPWQiNx8stLJ+BpXYNIIsvjvFHpI5tbCXB0ozxhv7g08R
TYc8Mp2QXQ8RPcXBpnEkEotCasfgSkBhe/F1toCUY3QE94Q9eoV+gkbYHHy2p4O58GK8YAZDUtRR
tYp0T9Xm0n68Ya6EiSllVeTE22WsE68VO5t699ONVaDX/2CzoTqakLFCqeX47w4BuIBO3b8O7BTB
2IqYwnE2Swgbb/m2tGXvOSrGFb2QwPrDyczzDAxg80VEZghIkqE6uOHzWTYQYb7u80/uwkDKKRza
dFMNnWCKDTVgC0FcBtoUhsRfkydhfFnhdvNx3gGooy/Bcw1zdZMu0yKRF7MtpdLHZi525OycuI6x
CtWCwUp7ouGQgOsObHuZs8IgiRSLa+AAGnLW4Gz+71AG+vVnasXgQcShdqO/OmbXZrFSvXDO9TTb
viS3fRQIBua66X3x3H7xHHsmrokmDaaClvE1yQpXfn22uHNXHaC/nxI+x793oRBr8FmAUegERMfV
K7MFpIcoH5buy7k1EOY1lgk3aOPKn9Z9mtpjUbUFJTj4hzYa48wJ/YnYzGTrw0JcBsUkYZq/jhWe
K+RI46uP9yhzsBqv3k447UFoCHhx/p0PYx2sufd/tCwniuG7phsl0CjUK7C7GoBhYSQaFb1NoyFt
qGskFDUgY74zM3iwv77z6rgAXBuwhQ+8hZriw1uM4p6LAi5odf2KKmraFu8ynCBl+HKf+EIOstuv
DiHZ4sV40UWrycyO6Xbj6+DJ1Ii4tYDC94oiY7/RWg6bbJf+blEVxW8N5oWqvHL21p/B5j7Uj2FY
R3930GQiKNnRGu6LGwlI4k1O8mUeMJlONywZIiBIR6/PHXj5qE/hEFY5Jl+rf9lyFrZHNjnod3pz
YlJtajtQ85VCKbOmlbKacUb1QOg2tyiypUcOl/BKofIE7MtxeCY2Q2Oh4ADcwK9xUDiApFZym1RT
F3a8XZRzHlHiWthqR5mu5hcWiRHdfAE2ge+okd2OqqspAEmZ/qZr6Egc7O1IQIWj1VU01X8Wgl5V
XIekJuYG2WNBSbxcBveTKAVAYojvvKGfDzAUgrJ8FhtXPebDQlTxDtKNV9dOSnqBZtjU1gvgB+Y3
AAqgo9TOpFZJMZJlQr2/0PywIE+hVnyqoX3VlV+m8N/p+Ud94Mao571pjmLGcd20fKDTHSbMfxvV
NDhSURYRTvrvJtbPxj3pCrrBSXYXJje4c7U0T4PSg1qER7OAywe4Nf/hwZNN3Mt//pkZibHyLFpb
wTHz6Lp6ZvWDueHXUY5ViCk2lcf3cjzeIu/Lkjh9sa8FWqFd8TtAWqUsLUP17k8BPjfPAEh3/Wx2
8HQn779foZsrjOTB440VLv9E/Hhh/wV/ATiLeaQFF7/cdbW6gzrQNva47fbOFRrYw7PRDyhT1fPq
aTWAFYmsndsfvXcs4tWAChQ02LkXeFdAD7f6fkDaPAmGigxEYCZwnRg5pPM9jaOLzdOoYPUOEZKf
VdmzshnyFhy4zApfnlHZfUb/WWtF824thp8iHM+kgsAn+PCBSWVMTVz9kV2PvXrUJcNF98SuXKp9
tfcpCaURxaNcvIJDEoYrYBkwnPUoEBt7yK10ljCiOkgzn56y3+pglVDbzkB/j72VNbd0Fdr8k0H9
jgBS+4ntaOGpMfMO5d0+JLygGUBiavvCJBEw278tax52+59F4gIp8sYoLw04a46b+0tDzjDSzO6E
sk9C9Mm/2lq9V0qR45d1gwu8eJ/AhfLTEBzNm/RIaAt7rsUDYSXJbB7ZQkQgrn47BEFxMvjdwZIG
o3gnMVtX3eOOBoHR+RuJqOv9hONd2HitDca5peHK438RR34VTOadjhNUlYK7i0R5pRP5ruIbaeca
vrH/snyV8tPZN+JPrFuKH9Uyc7CkY04lE8tM6EhnDVtj/gzgXQE8NoJpDoZkqE4Ri+HO6x2kDJgW
NmdIeMYfEJLxs302aqYByDoEeVR/aOKwGyqRNt7DZTiIvBdbKwwz3mxbCJ1SIPKpUd+E12c13/oB
jARSMJw3OZFiF+IN/L+JtnN+0jf6kxp65SWmUOVNNZB8NNkioLMW48Xsimy/TYXmPVcCJQG5hSCZ
8hEwY+lfA/3527Btc/1pq0+eyXbo8AI1kUB1yCFJtDRsphW5oYeiRoloq2fQOcIVnh5WySLyRYwy
zeBu7GnPonJW2XYTfQENbDYsyS9Ba7gyo6eE/ma/0Z8shXBy1YghWta1lxZcVunvYxnnhEPkE5+B
/6ANPIn+0FC6Efk5yxWtTTCkMnLGYX4qzap2F7iUfZbCc1V5d3fAQzA/WuAJWu+X34ZCZGtQQR0a
JKbsZhEHkLyCefaFqqpVRqteiDkMR26keuNmvWIlo3bq9G99V3v6rD0iGVmnhlYwmqjIKxDWbQhU
GFRjwQf51yGA9PIhOC9n9PVkLzIbv5dRESB8GNvnVZNfJ7D2tEJVyKp4xUZ3mml/vupffNFIaRCP
YHFUt3x2JeWZPqefo9TWbtp/zPvgiEpXxr+AyrJvWmsggjCkFu3506egcDMlLKM6zZwnmjs3X/Wp
oYs61fHvhS8TvbavwuzdjZMMw6cHF4gL43POG6uvg3cTMkg3XJtCF9iabEh7M7ZDBEhl8Cpg7F+n
OEwNmOp2SSM6d7TMPJqfHO67igZF7eg/5EJp+v+CTNy7OHQSQpA1So4r1hT4aptfBL0en93gPFYK
9BwM20EsQoTAUji+F3osD45yKFlLO7X8Xy+8biXXlsM3QeckI6wovo4ly3esfyS/SqF0WovzOGQV
rXwaT1PGa0mCEPBlhSWONQBAiYWRX9pXsAUd3H7Lnp2mQI+FYaJlaMYZCa1hUcEcI2FCmGYhGI6f
0eo7+qDkNnPe9xAjMptPKV9u3ahCbEM0zkQ7y8ksC442Vv78SeRA7cWbVgu7pgx1W5+21z/TQRXk
K3zqz5y1IFlnKCMHFSpEryPxK6mA7+Vy42BA7QaC61/yfNRndieEwTV1TxpahQDB3/7ICoJ5SuEH
25zQ1dgTet1/BxnELw95W04RJXLigdvYmbWvNJ2dnGlpuKw87Nfrmp+ik/tCzJFQKMRAeKWCAIol
A8S0xrhzeN1JKtQSnBXyGcxLJgAKEV0N0DrBNWDU+Xu+yT1iaHnEv9Ik0sffoRxloyG+kd4bhkwJ
R8nI+3AZBhfYkwhQ7m1wjuI7vw7qSjEA2MUAfWQbi+10FaBu6z6bvGCAPlsEwqGfjb6iHQ6MujxN
hJALJy0r19rmvxUkdVBg8vZVc28cYwDZhOaE9QKaytU7emhiJjOOd/i2SmJ+aqrk3mN6t/mOg/ge
B606wYGGetkzYygq4PQBGBo/i+B9VHYYTwT0e02HKU2XolMNV0rE/O5p0iMtQYQfSuVP4l7Q7SNo
V9A5LFsEncTwDxUwwtiUcMk6IIe9uRRz6mi6wyfVd9PshQWtrz3Unw4Okcm9XjVV9mdwxY/JkrrO
otRepitWDaT+FAeY0/jeCwS2VuNDSkw6VjHODhHIeg/ZOatge/9g/TchQcnMulEC32uUJl7MbINl
jPWB/XX6UPK+XCDCJVDcxcMgBvUznzXEGSVH9NidPqTVJRW+zDr6RFcWBL0q18DUq6+wNnkTQ0+X
1MJRrUJ98ax5jVjsU+B+Dmm6+vZ7NqGqtCO9DrldRNgcxG1HGGN53iO5mk5AT3j9DMWInFVLjQAv
wsKdiBKDV0BfdE0Brxl3yalZocAJadWizdewoMoNVmRZ0M5xim7R9qVlfkuxhOBaJUGmYrajDvg+
T0vG8WmeN3rUrpQTasEp+iHfFyHLxK23sn7M3zfrjlLIEIwNWn38kB6TiZGbE6GY2id544m/38Xq
ajm5RiYNEdkupeiIE+hSz21QXHp+T2dEIBh9pFEl/m+eMfZy/ILklhO1oRplliN/OuhjqmpktPSE
ZfVd9oiatY/TCeJKSoQR7bAO+tAAOG2WN0Mib7mADDJd8vV0Lcam3J6EgfPd2XPRcf4F2KlX6cDO
YJG5EpixSnp9ZtWkT6qtLkaoLvgryRIX2FF/MysKbivHVEEBMlLWoAkYL/Up7+Djoh82+KrVURzO
3sszrU841jqUxVhFxka4Mi8blbVQnYBY829e/1hFjpGezteifR9qJslFXqy9KGNzddJ0nr/CJ1KZ
oF/YPoI/jFxkG8urZoITiLnYMVojDIJf9E5619QjgsUz3NRC/PxI2m6LYxtvIVxQvZktib1lGbjm
Q0nkvq6OF1Xb2AU/BFykA3bxjDfivpFBW6kf/bAQa84GJdyK7hnEM5SR7mI4C9sPGZ1B5RlSP+//
x41uJf9PMQ8GxTX0PQWFKCtecLRLzRd9x0/m63pXMdC/DJCYCwaBglsGAUq6HEpzlOKPNOOJTLLB
DrZXYUCV6Crf5RZbqKk2uiJfLrJYUAvQ839GyQznSWI6Q6kHbUHg5alAhq68NkniSR0qIMVgiJCc
s+zBZ2Ju48A713JZuTU9MSIkEzdYOkofyyJlnjR4t+if8Bb2LLLh8Jbe6AUWO/fSw7F3fXmnBMbY
BiKhIMhPia6dBvnX9lCloxaBSJMxN8EfNh3kh5S01CWUeHs7CZF6lxFO9ExmJaNNSZvSgssxxyYT
29uBH6BDYV6maKOEQEp+XetMpoqRDJQ8wJNZmGmTEGGYT/heCjt5vK6xnk1e/8zOhd/vhAZktm+r
evxiRDmlysAqvuNeUhU5VKL+jrIwYMruzrc6Fs0b6+B6E/cB0kCmaywWK/WODj4NtnGcOXwSfR4r
no3+4XRMpHJ8i44QjGXyUr3YFeSVbvUm0jLX/Jd2HyLh7ZUgcgv/7rV0l29EhT+InHLvIoemdFWJ
Zs9D2Z89vb3/2wpTI4/iFIzyIuu51Ozc1e2MW6khawR7R3RHgZWqOrnE1Sy1nfnx1kZWAy9Tv+6w
LdnhaiVz56OJGXG2fRUUQD3zsX55eO4qIDPxmHCqNxROaz3tnTNl6pEK+tRAV/IbUtpxJC3q1YuR
okkUI9snqXOLeuuJd7bmr8qacZPbDmlL6WAtoc6uu3brP3x400Xyljp8mukMjQcQbElMKHfZ+AwN
LzKPAB2sHpgoS7uQ/GB6yBoIS4jPVa4ojGcsMkw1Tx624wrjJol1IqaNfd6XYZogCSUN4nKGK6i/
sxTLenT27Mozv8gLJZ+f2MHn8N1pJ29yEYFaJqHU6mtFc3ORsQVZ520/faPlV9kuI9SfV+yAJkoF
P0q5BMhD0me6oo2qoyP+jFp61EKuX5ScahIrDhwoXLesfn0XFFeQamGvKZtIIXqJhp4yrt4DPnxK
vjbMyMj8OiH9u2XpX20FOydyECoegyv1devjqikbynDIBiiUNGyLtZ5yCPr42/3SA1JDhPy43twN
qCCv0ilPpDsnxtZdoDVTFyWzJKVPLGtEbkSD/o9RBy0MCtsgnmfxrKqnyi4RjLGCUekgfHVlTcsr
hd9QxH+kcFTyDOonN+GAvLpZfSrifsDqxb/ENlNEHgwq/N3hTBB3T5ags3EHNE+rugwDJ2JJSZsx
+VIQ4l+DeO6Us1FKsmsGZtxck1SlEPLkCkbMAg9NthyvQcfNMXXjSEzTLGgAX7MVNbIfGPr6IH23
Yr5JOWn+lksvTG20LpNn79wzyBArs+cf2l0trCXiu2G7ITVDYjsuJmECpH5hZBOwTCZaesP+ME6w
UOUcN+h55BPb9fXVw0EMlKkjno1vDSe745rywJoeebc53c21nwx3Nk1Nq/oDBC12lP0fZo8fgKlt
/N24wSREiX5huOH1lP6XfKZxIwdVkSO4/g0ohrCrKg+XFvoAvk0vbOBHnNyR9tfajYK3jqkBUVdp
12QtBcbvEwuFUckuwMsKGC67yuQa400rs1E7dzOEhmypJEM5skZlYuXHtoU00B5pD/xZRGiO9zZ2
T3HHkPfR05526NN/7qvI+479Fm0MembfQjCO4+AnK3Cufr06SUFrufccyePjNHJodEBPdPk6I5z7
ZkjM4j1xWjoXNYJL6kE4oi4btgC1tbc9LZrsn9dlP23VbymKHVfv/ZJwOeNN1lKQDWKwTRYoztbX
GTdqzNQmPyL6RLjCeECws8fKStedTV8mNI43ytFky6dqGPRv64snz1MPuvu2SP0eD38X3U7qOz2K
FihUyJtJfgzgdMWDjg7hdh+RSrOtX0+RTe1NGBsTESlnrZmRcUjgG8mXHb2J/cKsindt3iO/eA3A
wwtzc+ulziNvZF3zo3Hw61AyF61HvlM7EHZVMC/QuZm62mjOIPoqqrNnvq3+G0bgx8ugpivPo9sW
7sh2Caja0sHt2rrsmwqiisA4GI4DkDWrxGHJN3askn3BYCsx0VFT0MVsSF3caFJG/5I49NQsMSO0
RHerClwm4rcCR0BrIzmO2JHoNyF5jmtC4SwHHjuDDpvHmeSS+Iw5xoYCWSKpnyLtTtjLc8WRLlSP
ORN4aGK+KwA0bl+jz1bF8zkKglY9d39SckpIyKMtsSjFk4fuJqkR5xtja8JZQa4ssGrgQZuxxfv5
gzNISqzTNzfSpw6FnKU7k7mW3yQYBTLHMjfxnbUcr73aHHNf0LECB2JRlk+17WxlS28ZuQFk1f7t
DBNJcLIlHIpWZMyWU4POMEGYB7HjIASAQ89EBPjkWHPSxkEsWYsbGu4zV2RIZ1coEs/sXH23ttT+
y9Qnbp1LIS3i9jbYY3CQhZSLgB0BFvQbQI1/o+qP7MJ/LIXLf9ADLhi8c/P1MdnuE+azfu2IgNFw
0TGsFYdQQE7ic1NbnsObHfRQPehGnz8yrOedg9jSh8WAq3VkrMGNdTyVcyCfGbG3G0GR3IEYmL9z
JQEfuqFEoEF3itoJgJSX7J0+hxo9hkKJ4FbywuffO5Klfd2jO47qjw7wIj6ufoQxFwBUrA27ajyX
Zqp/ZYaTyXqKuATeV8UxQ30+xokymC5nGKWiU2NP2BjIL+t4NHtSBCq+lekk6Iwgr+WEURpTYjDF
sMDQoE34xOEGZelrM7TxEr8Ed0MWXbiPPhFKk/d+pX4/WIkOANZR39EWqeQKvK5NU0bhknwNWx59
FKZVxHkt5lIh6+qLoklNZVtV97aIKrBkdGwNoLM/kW6dFHuo6V8x4e08GKp7KmI1RDfgaiBuzvlH
q6MFd1iNe8wXBegPQ6meY9VfV3PhkMJloJmdpShMYdUes9Vi7JZzbL7zC5KU+3FlcXpeUfNwOXUF
sLYIA9sU7iMD/N64zAAvojGSTOk3wk9mGt2AVJjhKTDeYXp0bRMRVkV2ENG6nqNxAsONyFxEggX0
TlsLrQbL7uDM515K4TPALhdQIPlYrMQHEJxZAOfsCHvkCnOCzAU/VmiDlmRSAhp4pCnpw0Z6Jys3
frhH6vwL9q/3e5SpaupiXrP3U98rUCoWrxUZwn3RMrOBUdpEbg5AmjsLULpgnzAB1PnQ/vCFg6VZ
t/BC8HqhR+F9+Cif5bFueV3RNHJHRCU/BJWFczAycLJwnRaJIzPIgo0qn2WoprtG2KfEHUlv6Wyr
erytQeVyu6DXGpQlBOTI9u7CXId6v0IjFX1coy02mduNj/1gS/yIr7S+YZ5pGc8ZUi9RaVQunQHv
gmqFcvyC+zJrd5INUZZziQ73x86vQ/RPX5IIWL7jGuS9w6njcgLnMD/ouSDcCWzk+tZuCbiaekTi
pWSBxrsRXXqk5exRas2MI41k2F+oXXyus532flnw2WCUtud4rENxojI4HaTgWhGK9fJ1yuehvHmr
kOfquJESZYADPYuTdoombaf1qgvHGUcpSLPLzKts48qweIA1tGi//f+Glt1gIZ8N85KTCUNH+3FK
7olJUQOYGANT9uMhsPYhP5Y0otdbUlTSL5Qw16SEJzx9q+6SrkVMGQVPao8Z8yZJ+8JYRjrQ3fOh
bxSNctbWwfQMcAqZyOQTotFIYUfq1Bqi/th353A3AfGEfee5WRqvABucJiKX9gEfhT90ihI87Fq3
ZylhxsRM01sjGPssLcxDjbhHY6SzSixeJ19fzfTALCVHVaG6qZOuvQsA1P+VSPap2iCQ6J8hhwNb
LaC5SvXZgW09c9rcq7eZnsh7yNN66Lq/GhU1n8WktHHLLGPldBh3As04WRSf2x9rpMFeNbdwBFVv
1DNHKvJBGqHVoh86jFaj9FqzB1oKl4UNgaw4EqDC9VKvt+AWOscnkmzacCyH65RiZUck0N4Bi1S9
tYX23amS52TVqgzplICOlW+fzAyg/PVt4D+eAb2NNUesQkK63as94N05zhKo8unG4ik2gzR1M+uX
qsJWb8ZqbxlMqB0PEk/+UQ/2ZAIJa7Im8d8fAMnByJz1KTeI47KATYJRhu2jBM/qI5NyTXsCrc+k
L4Zbu5x3KtqxKEY1GrwbQQ0d4j3VExQI0kt+511St2PdI68udq1ATAwuFwzcm6Ve1V3tBEI9TDtW
W4sfG3bEwJNQn2JVjrss5hOii0PlRye9vWC8/47OJxD6MO143sjW56QszW5t+QIPU6cgpsQYcB25
0Il/equt2IubhSq6NGZaub0rq6JmAC2PZfPWCf9EiK8Vt5i6hxD5S1PFV3ve6PgUZos9vfuShtgJ
9ene6nOxLsnx6ON51gEfblzdgSUWfzhgFh+WwYZlej+diFb9tOe+KMylslXkGV289w2dSZsV1Y+w
D6EotOTdXUhokGaVWpUb9Fr31myNRR7/hGjsNB3+YzZHG9T0O9ERn0X8jUBBDxLeBI0Q4Dr7j/Fz
fTBOxVh4QCrmK5rJSjBcfQuA4+fO4nCB3qoxAjG3aoMHQqTMAX0cggjMFQ/shuEuQhMebND4ysVe
3CDOdXlUfRbiUylcnAfJP6Xkxg8aZjKWO39BF2kuOFMq4egjqf9P2G0Ot0E3ToxigjsIevuHC25R
gXoLiUOdYVPi3feNwzOcHhAFlKoJ1F/8jCi3OuW5xZCdY8SvEsN2RQu3s9BT6oMhVhT9oTfET6Y0
un2Ln2U1wYIFOtcGHyn9REFoLVfyp2EEopQ29TgLLCfIAs7oQLJe1ojCJ0AKu+n+dm4xHuAgY4pl
KrZbDfXAU6vvtuB4qTMqMJXcILL/aJsVjRb/jV4H8u5BvxL/f8MgvgtwsCCQvdsgfzz37B5h8LhX
NZrTZzGQWominLx+zyKDDoL72hnEb+vlprFm/aUcqUa24As+oRAY6fd4caEh2nZSpsCMSYIaO5XO
XfQn1k03pDklnvVMZSkdBbqRyPSZKNQF4VT2bYOQaWWFEK5vYQGc8Sdr9rWSMcgVgCOE2+RPbBoU
2CLM7zSy0uMPpc+AI781n5C5Ii39irDkrDbsNMZ3WyFg4go3OZJGTGvxdQGRREpqKGu0QB8aLr2f
aJG5i1u4oH4sMhTdjYR+loibDLdX/B4+r4IujBDZVHX3TEmLW89JRGg4gILppKUYOaZrJUneS6P0
EPrX5MAC/4I+j5VVL3XjeMn4BvcWHwb+yCzyw6BvULoX8ENu1oe+NrZOwKUppUpLtbV7PKwjml58
REmKhAtmfKcmDvJnhDukwouQdAsymwgLqItJ+rwpKXSKEg0FGxjma/fUQ/rfOcIKX0Ea22Ik5OSj
xN35sMt0poLIR4J1+I5hNodcgOPYKReRQpyubVcbTRZZg9e64pkbGeLomJJdfehMYaJVveEOkJaj
ECq7K86q+Dh38H+j8RKIJTUo4ZiOusogphTA4Ok4x6d3rV2QspTX2DBiUxplz8RpH0+fqCnSzxJZ
22km1yT3QlgU5WAVD1S9KI+d8xZ+iQVLNwa9ncQXDSOgONK3YLydArALxKlnHZ/dtqDWrOBHfkQg
1dbnm5+pjHMlDfhCYVWe4M/1q1x1vYY1R26CyGK/AesPWCIjM3ku5DGP0HBNsO7xxpPeBvxiPjRr
BX1fouBo7tqFMdpo++Xq9oaPwsNU+fujdSy81XlPHtNvacwBPKcAkOlf5iPXDepbhO3rZqZ6vA81
LWj6OxKzYu3oxKEyhlcHeOUIyWFYJseoSQQLnqB5fMPNkuM/nqg0/nJt9Jz7Kml3TnOxrm1+Dj1S
A6fL8vYTvSLHak67MooGEP8hT/Xe3dyCqQYcrtBiQDsx6GlvGauB3Bzmfll+WhRDHqWaMM7TYrbF
fCbhhvs3NA0glagLUtkpwXKsKgQHtpgOs90We2+sqdh+3mrQ19TKcaZDPw9ZQ+2LyI3qMSjQYSPD
vXDwaAfGFgLcqZ9poSO3DKzv8k3jTeJhM/AQhlcbn3sQgHFdLpD7wXroxkcf/lhl8FcQ1TSI1l/k
nPrMPLb0HIQJGOQgRvI+UZ0RxqyN5MmLl5I5skdXXAULhrAcUUwSiTRHnl1owkh8mR9VC6rqmqMX
O/XJPEjhj9aYZ8h7FcivOhgs/3f+O3vziN48DLzL8Lw6PSnjoVJafz0vtGk/fiUwXF/tvn4SsZI2
mQOTJuUgpEqvgmZ8/XVOPL7uX4o18SIU6Q7/VBEW1iNqJtWr3szVsG0b6srG1g98c9Dn+cY6i0Zj
dLg5Kid+5G4LQsu61wOF3hBuzuyyrbkwjEfhFAaVyehvWn7ej86xJspo9g/rcst0Zcv8yiUVSH7m
0I7A/mW2wjGR3eShx0JZR5DPpdvN0xVUl4p1xrxU/lyc1lDwiLZ+vIJYYgNvwEFob/oBr7ZV/qnX
yD2iuuP4ef4/Zt03CGA91iL8m7QXNgPTGpW/nQv7ubO6mHVcb18cBMmMau7spJIDSZJep2KEj5/2
T0/jw11hhFjRKGBF8cXjZk71tZgncAyCQdK9JQyLMNDgCWSSvA3mnBxKP3RNpjYe0FjfR8jH/oGT
qVK0xJgqeWGNXj6MbIm79IH673zQLGlQvHbRJ2AFr4d3fQEw3JaC2kzzQo9F+uO6Frds/lLEyArx
dOGUbU07L1sxkMBUT3WNgVoW5Tq+TS0DSWo5z+XGawrg/gicSCecZPV0k92vVa96Cl3oGdFlWegv
PyEHsgBUC1xQSfhnKjHePHIu/gQPMguHziRGQ3w0U0J5ZKk3UKJsk7WN0pn+Dluuu5OMzmL4pl5R
yJpFTMvxfYyMmHsbjgjfe8aOUqBfmIM2ezd1PccqSB7n0Qn8CC5iaNZf3b1QMOjyyqzZ/y7EwJmj
byyBcOgi49l0sgLH4NI585pww9J6y4KpksU/RJAui+M9zGk2/XfT86bEdPyJnqqiFC4ZWOcHF/Yn
g/HZLwRw6QLwOVU3g8C9gT6AUrhBKNpWkIL7nUS9dYUAwKxWlBvpV4lXI8MMOZb+aGvl2rwUWheF
/dq3B/xBJpxXyK6yFwLa1Gquw8M7CVmA0NOV5VZ0hWh4VuFmo0OOPPqJujtrTUxk6YHSRtIIZ4ze
Xz9GZUeGyFa+R+CluJuK93eLOoa9ZUDh9gOakxNbFnqJYvUxtjx9bjcZleJx0W6dCP8nD3RpRabB
aomsKlSAncUU9jZLioEoU1aqAmLUOiBqxYRggBPRSq3ItPLiQfJtst7vyVMQa3ByIv8XLsH2651w
QGJM8+Bn/Vccz31IYNTiWQtDhH/95Bw4JBf3yw9VTwMmqoKfTR47t3g3WhCn3Bu4BouZqcifOkY+
48OPAjvUZvE4HMbWqreg12xlX0G6agNkGw7bdc2GaAXcTUUcBCjhIr6VtRbDll8hFqRpr07G+yn0
oPSnlHPZqkVpdt096JUIGJzF0Cbee8s7aU3gnA2Gc9Wj6m0AchCuG12+JNmwJh7VOOh8pnJdHj6w
tkCBGO7H/dcxZLiewOhUrQ6v/zzTPVM/ShsR5OB4EF+8qLUVKUncujD/7i8nb1VNcme6QL4/iywv
Hg0ifMiM62IByAkPSed+Q0M40/yUKKjA44uaROu/hEa/nOG4iBrNj1rCnHB4RtOFIpVk3L6JCO0x
orZgfR2OUFHRHXoX55C4RKdPMhezrNuTHJE6oDphuyfr5HKywKCEvfmk7am+AsNUVlZRPYxBEV+n
A0tl1TXXTI7dnQAxlLBRD5X9Ugj4nhPw9aCrqPRunNqqgAFsaPdbksbby5sET/X9mLDEmRBuXpuo
f5cmzKGwAb7CDbIMAQ2pMuKQx7zqUsNQTPqGWY76BRRE1YJqGoOHZ0kb5BhuATFxlG5ahHXdcpWs
obw0f6iFeYAEgAgKAW3I71oKzb/EqS72cK3Vlx0/y9wxKrHMEjYbC0fp0Bv3gIx1xzs4mTbLDxPG
6iwuc69d4ZHgabvR4kBbQ3sRXmEfdVjYPWc8bvKwIcDmvA4JxUj29qVSFtposVZkdOthunj9ggOy
rHCpFaol8KQ31ytGy33POmTO61TqtCsn4OWV1gqT9g8iNk44i6piwI3UCnfxxmrSssyGM8JNXOsy
1KEH4tuLO/w8Am9+OT1HOvfBio5gm8OB5U/l/Bd9fiymOeaTAsKK7Qrm6wdpES7ugxt10Yimy9do
2WevAIK6otUr+sECinD5gtqqmhFjHKbcB88W4wZntTZF3+XPcyOjN9YfV65OLbmKvrEcmJF3yfDE
Gw1Tn+J/RRp1Qbk8xvkLTwo2G7c3Vvv9/tQp3HC4dd0++b7RMZ170WTXd33PyX+2OQu/YlFEU5TT
hL5r37y6b9Y8NRxMWnZE723o7VG6PjHj3g3lj2of+Jlr1YxsykKojbyHaao+faY3xDEe+rXoki5N
nykLFmwgunNdmVsBQHPQsylBkZ2D5amSQE8ftB0VV9Cf06mUrQXf47/p6APSyG+VPydtbqQEN1g6
SDQ4rSFQLLR30yC0Z9U4zVwiZzUkZ+TRtCP+xW9MO4Hku61l/xO11hlkNiG0Miaf9GxGIu0YvVX6
f0aOqWqRxQYZrIPFP1B4PFj8VX/MxWilyZyPfWXR2L+QNf2WhyCZ4r4U9htLqF2Om6lYSTsRqO6n
FnE1BdZWjdoGaG1WDfxCxnrGEWxBUdLR+7MZaO2AvBhp3gPNkVIm1Dm4n6DGOdcgjSd5dWYBykQt
jm238CYE95AzcQgaCH1trghDAxnKaSUcvUzmqDbpgTXlDWDk+TY9TwMRG0vPnf1s1OSyFujQni+u
SI4DcmhHiY3jOTYltdjEbQjqBUsZY6TUqmcPOxluZtZLsfDkcGPlqk46czPbeaepl68KetVTjnyP
Rzd+XD2vyfkiUsHmpKOR8NcK16ZnvfX5SsREN2HTe/fYbBWxDHvJch2E3rx5KSKphdiyp9aOJnPX
nWCbDXu9kyJT7BV1N/aOF1szkE8LYLtX0re2YkwIU8kAltIXTEp1mCiBkmYFvFShFX/d5sB8qTsY
0OmFf0TqmdMN3KVkW6qSrocJ4qCZNjZqQH22L8t8wIcH4ZFP+1m7EIJ3ghEAXk4gMjUmi9wgIPv1
6RtaZnG2o0TnNlyDA2ogjVE8GW3J+693f5TJ84eR7nV+q/QiMo02GlJPJB9KAM+u1E65zVwyHoLN
E94Dwmg+Om6qnAi1CPfz9Db0hE3bgeOPO2aSh39dQLLHH7iddh5sFy53Loee/uaBsEbOjR86IG1U
kIHj6EiMq8PRI7yX++nAwefVWQ02SUSQcv8usvujk3Y4OfpoC7pwG5Jpou79azWsx8B43wlyz55t
h5smSBS2gtsh4gBv/RyuHq01nl+iSW7LgNbrLNICeU/03GVoBwaYMX0+Q+DeTN8IECeWfxE53eW4
CnJaBMoFxDiP/nWxCHV0sFRAvNfkYM6iC76yH2S7siLeHc45DLP+oS4ntIBo6zWGNpDw3yYzkw0a
Nf/m6HhBoupktlp5TZv37993yijQpeg6uk1axJDya9Yc7V2QYkYiDK9vjc6HtWF3hgf5OPo4opiG
1tgMmyK0BOGE9EeUuYTrHuppbRVuGz0xqYgihjxaxj2yxTOkZ4SQk7eGFxp4bhFO82FHJN+Mlupv
8VW2ZdJ8BPNC7iTVC/ITWbHUiDYBrMcwBiP+2MkjWye5oCegt+4HmozGora7f7uzHfKgWCPkMXDP
M37VNqvIddzZ9u5l8ATwoF5T1WYduBEDIZe1cba7cvN2iqrtISry/SpfI1dYqjj5p1wg5K5uz6+h
5rjZEs6E84/e2vQRbhGB4rRXhvGNuj5mJJ8Fjduokrp5DolSQTQydjB7vNONMyh2TvtzaoI3WwTp
ZTprYOuwbB8vcGUbLja0tsTsExWLCcPrXr9Gf4hRgJmfrzAReofRqlhnZp7DV2UfWdc6qk5gDOlP
Ufejh8w9Xn6P7P94rdea2UF/+YJlw4JrhXWfO2xtwkvVknYjlibIBhDo3AKwqvvHO5mSZDqyinqU
qb8kf7vJlGjrM/rnlhXIhQiNuSbw1GVct8ldavbE5HPTao8cnOse/vEcRbuT2UtCEs6q62Tgx+wf
SxhTIg/nO/GIqO2d9jpGJXFCm4TTP1j06vLQx3mdROh60lXIod1l2aXggEzH7lYIFdtMugDuz++e
1lz2r2gRizOHF+uJy2Hqyzhht7PPdVX77OXSKmvlWwxL02kz73yMhGLsdjsKqJMtXD2muZq/4a9k
U92pRy4SdRDOWpLN5QL674QuTLHq/YzNTeJHYTgMB88USHLMsRPiwzE2tVmuEdgxTjvhSHxlySlM
dLU/vRQcZpbFu70VKeBsmoZWqnP3dKttcaV52Iy6pFLG3l1ci8ETqbOF4b7A7nd79/rq7M8TsSwB
lI0BW6mo/l2hK+Eu2CGh0+lrX4PeYjfiP5PVxrj8mxImfJq0+6Rox2IUd9fPz4SZ3DfaouTjrQtx
YG0M3LUVQiMTzEIRuYehnUOjMoVBvotRqtCsskPp4HeYUxtUQjkNE0H3RENvEyEoIqu79aNvUdGB
ZB4LGP1IWiIqw0KGmgtdxC4ZUI0vjsBuIJjGdKuJWxfqqTfncuobwpNVRzsj/SZytLqenktxoQxK
qC8M4z2+xOJrQTo17OsAlPP4r0fRnhm5B5Ur4mcHDIBhcTbeOaCS8Pd2MpXtGvZIQeubNVMQBMbj
V33esYWXK2mOhWoPCYf6bUt767leF15N6f7V1gIxkzotsa+wPLbQyfcHqeB2yWLf+3iyZJee/QDz
92oRMrpV8DxIR9I3mvIsQDACUKmnsVQJEZM1Udb/nd3qQ8d+c+HzAvpnIo8e0XY9F2h8+vE+gG5a
ebkfYtEWoLYRXfipgiPVhaYpIsZj2ypg8MYrbYXs7lYJlwp2iitCP5+Niu9GLYEg0+FHIWnRMObK
5QL4Y5WDO1EuidMY2KjCuYGh8EVC80rX1XFwsN60MSERo1kER7dP60hJQZOqIQMKnq0vfc/6VMga
ZKPowbqR6OCRfQwtAr9IM2RHHWDmtaoIercIOuRvmqPxQv437AJ3aUBT08Lc52fhSBGO6UDz8AvA
TUDONMVwx82o1yqJH9VFlb2Kpq1HNFzIW0gD3eebPIxfWft4u9p1FdV7RmFU+5pUEqmStv3YA/T5
ROxu6gLzuTcykz14LVeR4G5XBhUqPqLQ0dUVFjc5u+2lUsW7qrvqO5VluvC08u6Y2oPD/dbZvYue
c8690jUpBZFncP95kp+xUNmBAbZsp+zZiPCrhhzsgJHuU6gboWJ+l7PiUZccWgLbPKWy/5gFK4X2
ttsopo6jJEoG5aW7yYoFCMRiUCZmARymQr5t9+P2zs17iOJppm/uLfUDLCPorcHANCoVf2gtNDyV
S29wf1oNjdMVi7Q4BtPwuZs9gQRaOcqrW4ulYxOpgOCnUVbSkiWjR//eQHPg1O5FgXT8z2tIzmdB
LWExp0tmgKBbIWJZcNWOb/Uu+mXfZIZZiQlcJyQIuy35vbfxrxYeVh4XWuhLbTYicc6RVNMeFVMr
3/9T2U790bNF3f0xbYBCjg6363xVQ4XqBj2vpvw1T+F3D2n49AyWwwzO4bIdjeO3xdba/Uj2EAsq
cCuwlylId4kcEHcRYcOmHWavBTaenMI3bJHfyusP2c62jFaaqITzxsCVWIPTtseuirSfBEGpG2Kv
YnTK9AKhb0o2mg7hrJX+XN/6i2MMNKNP/fv3XG0KvCQR6Hpur9bUgnUNKJ4BANAMLXxLz1OCgqM8
WYhFlHf3uaQLzpMIcN/IeELV6dtJ7CkF4BdCJh9RpX00BDqR7jbuJVWOBXmMSpGto/USsogVFXZg
Q/MXEVbh3e8tuhQ5AK194bO58qlKd/g1XMzQQUNSDAJNCbaVvzyBKobj7ogpubnMNoDumlzLvXPf
+ISc3bPLudiXDP5xdwE8/8gWPRqcs/aHMKiUPVOoRRGpDkd2Qzo79lIpS+JBDmot6UBlxKWGPTjh
lhjD9Rblq7odlC27vr3luBBjyWKEvUIZatZH+XxQarUKBIFHdZEVdzt4nJFwZoPlmSj49XbD0mr2
pOfGmZ2khBXTpG6Cy9HdBZnV7X8rQ7QjIEzMKgIxjqpwlv4grRi6GG5FIqN1oMn7JTAFWgdvpfzo
Ex6zL74aJhx8vd0Osg9SXcpkuTlhi9XJC9fPhlrPM1kd7XP15Rh+JhNTsHx3URCn5K/Uh6Zp6HIL
jBOnTedTCF0szO3D/VGlHjRetswELZNKvYFp+rdDMy6D2FhnrDs5ed7sUrWbo3vmLUK16nEIBrYi
q+5C8fzRnseYo4GAdrKheQqGHTigZUd80qLA31o69sFdWsil2UQqgsF9Qyqe7C6P66UUjBAM/e4q
Zc9hpdK1W4KWZQzB5+zzFsPyAKRXh+BbGVFe6FL3D6y3MMGn+DxJOtqBDivASEswNrVszUWvIQaz
v84dRBoApXTdT2h7ILFDKUDVhtl6M6/beh/loBtqvs7FVOTu5J/bdYaMT7ZISL3LLvrHbUfqdLeA
8ZB8fPoubmua966xFVeIIFV7QQ9Hn9Kgq2PR/bhdmB2m9+Jqm7WPR5y/eDlGb7Y+2IR6GbHo4MvA
hmml7x7Cg6M4jrAhfQQ4VDDy4U7thskLEAwmn+ptbvMQpHdDbM2P6xyYZnO/gryi87NVwafrLObA
gqvdVEN+cBfVxwIqLh9Odr6miRSktnfFjU8BZEiWSGSMeBNKDUQrysbqTnY60jW4KLMrI/POB3Mg
M7bJ3thxXIbR+KsF2hCuQ0YOPQPswN/E3kbBJh8cZ3yiHvbNStCoiNmHqbgzDI0LBgFMptFnqfj2
0y8NhXpdbK7SOvqjKy6YO9DQRmKXr9/HSYcpc5owIUlv+iAGVxtgc9nqheR4nMnlNn8uu+UunQ/U
F/FWd6d5Zgme6lkcWeXGsMx0kzyXHzolTyotT5OpLm4/SPspHwimkHAcnzYI4Tp01b67mRooZ1vG
JQsk88o94eNmSsF81chU927Zmm6cxlrlX9Vk2syrn1xvKY2uIVdz9/0qDwrC7zZoHmpwBRsxHfrI
Z8DrjPbnz9F3oZSl1E9ScMcd9K2MXpaATt7eRGpKlzVE8EhlrKqSwbmGvkN/xj40dpG54koWZMGW
YHU1W1hvy7SvA0a5B+NdBRlFxvHJ2tw5YoB7WQ3odbLlP1vmjr2CrisrU0sHQn7AjC6dwDVtkZLR
QZsbPazXt3YCMKRzy3l01pC36ZnYmRNAv8l4zBR2FyR9TsM5n57vG9US/59qGjgVYrPJzIA6pqnk
98499jViH7OJetrA5u1POIKGos8OtO5bETS6V19n/4YGur8CQS8VVNer5d8CyTcDtm96XakLcRzD
2CqxAF6NMetvw72gJv/aWhhz+bDXo0F4bFxEbYZ3+dEG4idcJN92897BOMcFx+OINMrURL1dCphu
7kRuJp5xZ83hRnOzuEDiXl9Dsx+2JSzOJxcspYVlaFKAcT01Z/+8/RarPbRi5yHWdPbQ8/TC+CPW
E/+UuvKg2naEMbFBNIxua83oxhmNTgcUwEN6AGo9l69rINNa2UD1W1wwbfeU0o03m5g5eTCZqRON
kWrk6iCIWmg1Scnkf6tXdNUgsAdZdiJh8buNkYBd9oa45UML9gYmk4xQXoRCAkbLSEd1GoBrTetF
qEsUKaV6xy1eaEIDwTj6cjSHGPHqMhSu54HZjJPAjCOW9F2fMU6dTzL6LeNsx7a1NlU/N1WHxDxT
lAC3RMilkjW58sIi967NQE1Un4c5KBJIXbKKFcMBStxX4Sd/8wg2ytK4dD17QcKiOrZhreOoTKer
VSpP9JhzvGKtHBfIIcle/OWOK7CtNJX6va0vWbXFPJHJ4Jx1JICCUtDs3fjTjdGEu51NA6lXTrBw
L2IpWph1mvQkY1tq7jVOCHpRqNS94+Yhl5RvEbFc3u91D4aEiyVvPsgQISb9QxylKBID/qM5l+Ga
A8rLF0nR5LQf1ooV9DIZDI1Xs8P0RTdYeKaIr2VFrwWFJx/hdNUkNNm4ll5/ukiber1CTbbaEXSp
W4MveCeLRwiAg0Ej0KXP7l1uPKSSfxpjl1m5mB7HWd+WcdkQlkwV2K3HY5h6VJLM16OAZxMmG4MZ
uBv53C/Yi27zYnWqEQquzCgSbTS2XOVkktiQDTWFJb5SqEiAPPubOwzVMbIYbuWmbj1LLa3BS34c
nUDrhHESuUsf55tTF8WBc7rZTKwXjDOo5hoUOqg+Ti/lnrUQzM4cRZXoP6cydmmzBJumABC70SEF
EQDsvJXL8jV878s+YCqaBWt3I15xhJognLgfVq49/fV1LawmaR9q+e8JB0uAlPjhyW9Vy0Bzc8X7
hrO6Bqhde6jLrxk3L5wGzfocz9GjFYUQnQEfHY4okOOedAeNtIHZrCE+ptcdyvXklSB8U6AEUgKf
pS808q44/HKSA0cACrq7wCujkk6RFB7QKiNuPzY+E20AREzYOzEAXpNRq8ogsyv/Ys55Q61FdYid
Eiz8cdMQ/KoPI5DMFgI9OxIBVhcGT0LS5afoqeSrK5dAzh0qNTG6bcWsYjVJLU4HHPnlHMt4Sgaz
NMYQ4TqNMwJOF3CC3624unQTUaK36RT//ZRB7VPxt2Tw3Gx+93PyAdU9+6zfmZiFZgyLnNe+znYX
mSev8OpPb2ZtGjdNGLK0LOcJ9FGkSjqVC6y+ur1nDnz6nngHhA8DxvG+sxfV0tUR4jhv2aCnXdaz
N8D3rfBc3APhVdlxhJeueiTVToZPNSWJfVjElxxmVeEJN3J6yGPicy3ZZTHu4IqvCn6O1GcJSa1S
VzQcRQ+HsEArysnlw0nz143rVa5l/T8fLNbANj7Mp0QGA14+WuOcM1hNB6mU1WtPgWq2kq0E5yRw
IbJQmYNealTwHG2FlezNwgFZhT0LMMD9hQDjFdHFLCEtGvneQ3RxZ+8O3eXMk2n1C2Hf+1aFGNY1
7HBQb2xKm1v+l1kbAa9nxLUFxERbvlbzZonKT8zvgaEi4GLOZW1oZ44s7tgScmT80BzO1RZOpZCk
ebf7mp52QvoXTh3Zm5erBAXsTGIUrh/moWtm2t4gqkEpgZubTW337QF37aF/+0r24U/sxclOI0AR
pH1EMfLf8xwr+y9tgcJ9NcXtDvPaoCV/vKLqwyaMW5Eo5Y6OPqz25wcOEVDoqC14gtebGy3xksF2
7Ab2jvdFjyfSWW/H/91T2+S2RmdcF7wAQP+e0ECPTM3UBDGkcDogA9KWZdHsPnE7209MeNnVWJRP
QnaNE7xiwjIW3uBsDZXJMWfN70T50G3Gag/VWFEpW6BxJIOpoUY1sGY3dpj/DCuBSv4NnLIziKUp
i81iOc7FlxRA+fTSv8UIbr09j4+auuHqqp5omnTvW5xkqzptODfJogts+sYWdnsESYLVkdvblB+z
rm6ME27VjL5iY1QDTPbKKTjyS+iJMduBQi5MOjnfQBZcYeC3GAmZLhLmePsAEg/7rUJUc0eiH2PQ
KHFFll/SJyox4LHDIDlqcNLHpMgopotOSa8jVJEuOXIc2yUNGVqVqOXMU6BlsaOwpOzwSrwxH+m2
Y5grZm1N2v1TAs6e+dVR2qgLJbZ75zOp1UkounSvZyviYJ9R+ZAAIA/j5HD6TvXTHLMcAjMwre3I
Q0ui02Hs+EOMgjxsK4gaWGu23M7iBcKyZZ/iN6XcfoLMM7zsh3dx2Y+YpGLFayvsdveNORpfPZ8U
Ut/LUEiG4AhC62Jt/sJxOP8fa/vcDeyvJemKWzp9GnmCsJrlBAWKEnee5DGZkVK4kZF8jLkB0wxH
IcsyXVLI1K/rOuHv5hP0qK3/Dz2ZWFI3rZCjGtgQyjHJXoKGJPjEDiHurGZ4OST+45IjFBc/5obV
LhobCjBzR3djoK/oB2f9oy3eZTW5k6DsClrVBPBhE3gh+Q0i4Lc7dcy6d9slUS6oGF5iV6QRUBl6
+BnpjwC7XQ+Ht3Tut5UN4yz5gRiD9UWi4vqTuGhDr3kCJesTC1t/UZF/rTV7wU1FALndC9YCgLF8
dCoTCORv2iVs7ZsYxTtr69YK1tu0bWxhO2w3lBFcUnCfwSz1lrH5Mg5XTzGVMh+VCUYChv95ffeG
2gmLomF07XF0AHa1IMaeJr5gYwlMDxPpZZhRxf2LFXDY1vO8cbdugOePidfcL4QIZx82rHE9ze/o
fpjdBY2HCPgvqWKOja760N2nQbTKc0lGdxvXRgf/LlzdgEO8ah64QpprvS+cuuTE34Z9hOwm/hsb
Ju8gNko5J8n3kWIwfJKDD7Hya3zAfrRNztZwz1wWGIhldRzlVVtyJEhkrv7R3UYD09Vs439zCjp1
DgLHJrqsd4db9LRmUSmU+XJqxW79m0gFB7OQstssCq2Q62rIyHpjQAJ8BPexGa+YcOOqLZTxu/4A
+XF4cKN606HIG3qNitp907JifSLZPEEeP3eIPgIK/qvGe3wwqLl7VajUnwcXafmrCxZzISqlw33G
0fxLrQaQ98skpbotojsN961Ou5Zn5i/z8wBUnQH8cM/lg/Efhpiqg4JIRj4g9iNFAbCxU/D97M7M
rgX4EMj1JQsscPxV8nJEqc5acn1Ub3MRvv2r21iZ7HfFem8zlYIxGKH8iqWSehtWt83FSOAlQ/8t
q25HuoSe3wLZzaak5sXBwmnUs1AAalDTBTXkMcY59YiS3a2aRBplVBhUyicM12TYw7Ztn1GllCLn
KQKsqTM4ixucx/wJxwwzfYBOYkaVj7nwDkidhTBA1pJKAtqCoaUk9TjrkSZ1lXpLSeD6WYGKjAhV
jrspcuLX19D/8doAKqGkK0+pKzw1Dpv3rBVNZHorqWC33n8eEbvvrng5FIEX/plrRxyNl66q2pgu
DsbzVn6eeQc+pD0vxUyhdKIbl24hULHkUkGQWlKzwqx+SW/nyjom5bdOImaRMBL76bQ+9mmVYypn
ffoxu2RwZtLX8Sdq63Dikhy90Y1PHN8cUZ9VeUZ12x9PfXBtCEDq+ViY7qBuTln2By7cHW7avtCA
OYKSwJLqdouspVZzSLDK/T6541wtDqaVAatf6oXF0YiMIw0C2TubxF8uH2fKwN/hYjteg73p21J2
aO4fSlLw49ESLN/d3v3IcFPdOcY+8A4aXc0E7C0vyNqYnZa21rKSM+a/B7m7wLiZM2f65Cr/eGS9
e9DVx+WRFtqpUXk0nu2048dct+gImooKGr0alG7ESjUAdWlBMUS7ox+M7Fh/d1guyv7mmNY4kpi9
+C/Xx2tPEeHuwikjtsCAmly+RxvylMSken19ba52e+ruvvIcWZlBjTbgo9Ibc7I9+HfDfOj1DpWV
r6FYUkRqO2oEHJjTCCZw7EcsphtVxx1VGvc0+6FaBuUpW1fgB6Bv1XCO2OyO+PqIDd9Vw12+d5b2
zJrMi8R+9BUjt3pZLzpsPdD/7d0wtfL57cik760wi0YC/SWFz/Y8Tx9cx9GZR5zGR3XB14BO9xAL
7sYyseRJTgXSP4O5yIh2swnrsEUpl4LlP8iESEeSRk8MgccJNzzpHfPzQxDsQn68tdToGpGuxm2o
Qq6LJc6JduxIzqcM5driS/5Z1tPfp5ENZbg+i6XQSUuwPWagx42Tv0SpIHNImezq3ewchCyKZlbs
jaBJJRfG9kHFj3YB7pQVTChlBkvqJUnYNKphtaJx4x6kVF8vF+5DV2TFzXJH6Bkd+yDhG7wE7ii1
fgAxsYU0Xs4nZPB7I+eNCcn0SLh5NBC6UjGf2oDjD3JUvaJs9antUgHoHhLtIw1geIqwpCmlnHIJ
YYQ6vI0Ukq/cR+3In6KWSY3pfoCoRuZZ7RAphZl7lzhZYhoirOGwpsI4jB/oW/lzfWyzZroHeAlo
EbE7HibHp+eNUy0uKgc2LkgnKxgLXm/hNnw1KEOeJ1BkvKLpacVw8+9Qei8Lha677ylXv13gaPmj
fpMmUtS+r5745x+o2UrW+fabSyLWtLCywQKa/eZ7E09XurviqEN60Qr8yENv2+yWwZnUqNeWJJkh
mvWgIrpTfkt5noWN7/lGw0amGIrkbgsN3kJHgotPWwmwwaYIfdu9iyzLDPpyr52WVV41ZUSzeBdY
2QltogagBXs2Lhm41b0Q6ruwgogx3+FUTIHH4WX/22Qb0c2RdtLDZJUyoD9a1PDpw6pgwe8DKzr0
Pkzueep8t2vcLcFej5KQRjjKgZcr1dh5YZyHGwazXGsZcCYGVdE04CnTnFQVZqMQ7BXSSQn3hxCH
GPTFmL96n7J3KZ+mJ4LYmH8BGF90PkCY7FYcgBB2BJCQDg0ErLL0m0lXfZkFSWLqSGvOkX5D2lgR
QeQ7fHqH1lPQpJuXJ86CYLcUb3EVMG2wByAIhsC8JxlVfzCYdsvEHnI8b9xUyK42vRCZV3HsLpTw
9a/qM2vilEdj7Wiw5/K+JuX6loWnI8WF1jwMx58VmI+EF9qvMH1VoH7qDYt40oIh7R/a9U48OPAc
8iO3wgWdC26fVCVduKuaFMkkBpf+W8JuKIFMh3U5bZhxSs6dAHt8cUuUhsePBKZnBQnRkzQap7Ct
6mcAgF3JW8jTDbEngECcbl0ycssW1e7fQ+wC/0Mgq+b92pYpzcctK1f5nQ9DSVl0rUIrUQHzB9Xq
KvynmngLjxEaCutEfp5diMSCWTLueuejZWFb/XInRNpn0xqHDo3iqUmYBPzD84YUoOZ7BBTEkEyC
sqQ2ss4ZUJAaduhZYfZCJk7X5M+5zDPJU8bFb/h4Lj+lqXw/8vD52mh0+BeDci7Z90sOjou8AWET
DFy7lgy4vgACJ5pLtbsXnltNdWgFiuCmjx0RejCEwgdEc7kLKIPy662rQOIaMLXGrbINzHC858DI
JkRlZ8HiJMlnjydWRbfTDrWmqap5Mm3HvMyr1mUZqzqFuMwmFA7RjWmcnTrLT/FagMPitfsW/Fhc
jQ2sTLg14ZrwEm8K2tVMSqkApLiglxEL2vmb1oh4pGA6+iUNUrGcoYCExizZVkvdJwdmn5kvc7ei
83gOZb6qia/gCjVTnYzL9OWs5lVCMJ/kDoVFoIC12jVBRbDGqvG/svrjqrsu1Lv/aRdSnSNp4AHi
6lev+24YYiml6hjtFp88hsiw2AmLCTyOsXuiQcQtABP27WXUhRZB5jqOFecIyusMsxFaVI4DRKw5
SbT53u/trgE7Hf4Rih5EyUtiJiCbfNQGcFHlQeL0G8VfCl4ey+89dWnjKzbHGZRT8Py+9aTQAAYN
vvjTj715KUfWpMmY3y29osmPI4rO1SlA3Uj6C8xt8MWPTU4Ey7nPj8p3pxMtshV9k7iCHyd5H6IL
+cwnVMH2g0jKYxcoQC6aMKX/7fVm9Y0HEyb4ugcBLlLKW85j/BskVRxHVhZivBIERmNV6DBqkcL5
/rw/vqlohd6y7LPRQv05UcmDU8NIP4BNugQlcifJL1Jz8StfplbSMNrsiW2lswDYpAKg8fiFpP0X
aEL7qGwbGTKvXn0pxI/GuNJ8o2OQIP/Vj3kiNbeRDOP4goTULEvU5gvYSCT4kZCqUFf/M7HEsLpp
5oCUUpr4riHBiPL1iVimE3rwMaZYipg+ku7uZZOFEPWByUECDzGo1BOEXKMQxeIbJ7ZLHaLF4XmT
wySDdl6LU1N8NsKCMQnxLF7Emizz8dKBM3lrAlHU5FjTVaMTlhrXnPQwsGtIlEjx7vtLbANr+2iQ
BLoAtzqbBWMxJTdqhhcfMVnBThK0zJ/6kpwzTroZAsqPBp0XMGeDzGFzkbX3W+wjvWJ3HXZkkk8G
kWAoavGzEGz8ZRgw+H1JnLLSEeh7aM6biYa/tMicB0ofuu4kN/+KdFxA6tvsIQplQdK2zrWzGceK
cQL8dExar26+nh338TG02hYg1sKTyYAP2D6RiLEkcmYStm42IuF+eawcnewMqpgGzgX4Y2eIOUCz
lTcaP0lcxiqMOo47lUcHuRNuUzz6jMO0l16PaDmXMOoY/VifZwEHosR1z4ttXWmUTttzLyS58hKS
XzdM40FHIJt0iCIykLpQcNxuf0iw0Ec6XKM+2dPiCeAWsPl9Z5qDMgYPqpQ4BBz0etqEboOpPOTV
j4+DqU/ufxxMMxMMRzZM2oZRqJVl34sNGQyCEMPpB45ayuW/2hNS3PWFONAhIO9Mfh8XfjLF5g21
ZswaCokyXeFzPBDxfL+vehjn1C6BCkBq1gNB5yYEq5jHUY2bIzi4TTn5XuIDPbrqy1NgsJVHJlx8
ObupGYTLbVsBWszzKoP1MwIQXc1uKXv6fj5bJ3Rsq6l7CVTKhLiitwxCORdj3L+xeQ+HI6ekkzDN
Gxi0Q/RuBgjmLxTRZ+kasNuyZy/dUN/ZfGLwtJaGQSI5Z+iDKOmDP+m4C/VHBJpXKJtsAJTjhAjR
LjJbe02q69muGcBu0dyBxmj09ANcFdWtdblmX0gJ3RDLZznYxpqs8hv/4LOSvc+R7DOcaatuuINn
vXQ0rO10S7x8YH6Q3QpigMO3QUOAda6oDVE296eOf3W1iyNsgOvymqhZL9P4IdCD4ZaP+4omDuad
R/goFKJ3uAjWhaAYW3O5aicJlVSZgJWA6pmwvJE5cgfSYm+ODmqdE4v2GTpvsu+t9zdcCdRpda6P
1bIQB/GMBSEAbO3kIP13z+FHvfLFXBA+SZZ6IVx16lnNP8eDq/1oB2VB/zEluBBbsc8jqZZAGFpq
/BwH8kwyj4uNyfY50/H1sYA/UhJBBvolJhQjQrdBEz0DkoRzOtZKENaR+B5dNfSN2n8Ih1xzH3wq
UP8gNqksD/xKg/0v/4g7zTaQaMDb4BdhiHI574KbxjWKXi/LrIGQr9VUDEaTw/KtVbeSj4o3JjZ9
B1ZPjuMdvPJPta3vLxhNwSB8bGhenfYwSpPXgmCaAAZlMZ4ATUUbfZwYLFz+v5mTGcdFZTzHGRuH
XnA1soprPAnh4Am0lRoPFfCqbogcqFez0in7Jjk1Afj4riYXy48eRaNofC6grYXHF6L/qTzgW4vu
DsdvXvd+w+Ztuw+R/A/hH4YDv0hQ7JMYJzTDCG8XF+PgIycXlLtD/kl3NrOW1wzRPCbwRErs8m9k
E6dNSIx6fDge5tUEsOwy/pPOoYcKXAnzQMCoOY0opSve5qsyCIK39K7rQDNg5xbDs9gNfm45xtNF
7T+yPHcyST66WEZHoU3+3NY8+uKnnC9duR6yZmGFErRK6PhpsRqqviZu2sl+KyGZC8e2fh5OiFru
cpCR5029ObgebMlNVpOV+vLnE+cn7v0q6z4vy03ZGp8aJ/5RgKtzpzVnFV0+FIS+fMM1ne29MZ2n
2N9WXuYe5h3kKGP5Kba2SV4vWZqzWbr3/gwHV39+7GlFi5iZMrcLrqFq9gLlBi8gQIpwa7ek9vXV
VI+BRgGGWqZ1MfPq2JGb3b040qOComZiUvd1BCNjL7xRL2yzG2a8V0aWYsOTZigk+NKcuDhQzwtl
kjkOpPw3ySmXAQtV7FSs/yWPqaUI4+hHbnexwuMOQVSw8fV2J/Ti+2Rjh82tnWO9CK1tTYRfpKEY
/GX8nBrFAaL0pA2co1JUJ5gd8XiBONSu7zjqMHPpdHOtKv8sHwlm9MkiJIhsJmQWc8amsEwYgc4g
pmMn/ZXCIO5lu9Ob67xss+EFDDBH+hncGUO14HXlI9fNloJhZCIWuTtBCuoCVg1QqIFEJmfAMhuK
XO/P8BFqsPuY/UkZH5+vieCzpz0bnH2AfHKSkC3bBpnCJgXs8i58pctnFBerzmwp63DeKCvGf1nf
YkaZJcAfEpyQ/8ysw3OGYZgh4XNnfHTRFle85StO6vn/9ivM7d9lV1nKrUPdvTgDxiZNnI7Tfxfs
w7V76e8yksNNmhlyW4lszn5j3tyZ4aK8C4d2I/olFaxuJtT4/+nJE4ekjT8d0+UlywC13ujiGA/s
sbwnGmrUQoACnq739af2QTWwWNmyFkYnfRanKgsHNExfpF85cdyznQL4NfhEireNe3PBHwHsnJTe
I2IQXOqK776iWeoSbcvlzWm0wWPX/sQpLCRC8tVRkfrHEMpt/2YfrDluzl80JmcIJA3Ozj45pgJ3
wvhdHB8jBSwRUx4m2Fvh7eNUebmJKqBidd9Y867qjY96n79aihbiflZgoVOPdwTwkRDomVjIMa+r
KWjK+6IwxYwfqq1kvbv1uYxTBCsvQs86NbprDGtTEpw8KT2PpyYGroJKHPeJJgkmArZx0Cq26fS1
uY/8v/Ju1fqvrQ/cyH4MLzlTvhF43dGWp325KGpcrwXK75Gb1+GTlewcEfAlIOq229R+liLNSxBl
R5j+wcb8mhyjxA4pEZPCY6JqgsvZEZMKH78itfhS497/Awe7mgbVZTzXCqXGhopWRM6Zucxb3Niz
W6TYEfve/UHaS7rvvLhqcZm94lispr4X19Ki365/6Bnbq22Bec8do/XViLFhDJRt3zcM7FhGNp3K
aGdWLYF8AtDmPAWVYsQI34pFWjlZBzoiabKLySzvQoQYN6DAkGkp1i+7QPNshHKaxC139hL1TmNi
f2yH85ygXHq41dQIXsSgW7J2DQoaGiGOHEyR1+qJV4pCpamMMsQ+GreNNx/5ottAx2tc32o2Mn9b
Di7bc6yV22L53rSB7l+hJDwfcqBjITcNDgNlae6MKbppcfaWeIB69uQjtged9HGicbZ9q8GgwxWi
6Z4GJqj4rHoj9CRW+opLV0PuXEM3y8ziimlY7np/lkNcRYPsQwWMC3K1BT+DvHQ7oGPdj7ViXRWQ
Yh1dXmkRjzg4MDJqXobWcAvCTE6PBqXK8s5rnEL/UWE3dceqOVhjr5uqBclgG8z+CTnYLhM1O/Ho
ItCT3KSZAi8X3hiFzGIp4JXzl7iKXgP5ql8CZC91UcMSVwP0scgQeB4oRO1ne9uzsiXH+exwelzC
NVW7OJvgsaEBiiEEvXtsSkhXlWtrU3IrXONRiH4HR3JWfTUg1zDLYmnN0kCp5h5hW1uIjsjCBgbI
6pJuoAwWQ0imXxSoipVT8w/AafCv+BqXkQqS22fJUq66nrgD+BLl4plKkAmpE9TC+wu2kPszZxvL
XdxlaoZ7bBGrEvD8k2wmGpXL3LiXeWQ/Jsr+T/+sGoTha1WdzL3kGHglwVbgPv3xUbs+aH28bmfr
GHHeTl5Jwd1gImCYdPCG+sLPrExhmkGk/tBgLj2jei4emb0r7tVqhQVseUWDh37cPuP1n5bnL5te
wCaJIOPL2c+z5ddv0uc/HCSZG+s9ilHO+C34dI7DT/rWcoWNhy7/0QWJxqrfuSZ6PMMafjxdj74r
JMk8GF7z2e0EtIpjyIOxVF6niif1N0V2MiGbEOWrvmcFupnlj4vnyj0fHOzBr8ulAlNf4xyli5ov
pTBVlApmy7hQeQUiHmIm7D8zlCXgXF70femieRvwS0iyr0WqyajTLEUxTVzFLaXlOX4uHvpOz8oR
cyX//lFQYiwWdiel4WP68KDdzxxF986oUq3S38nQXaZF3rEV/VP6BJL9lLSu2YBcOEaqi999+XYu
ACwBpZEyGdIfX9xfDkSOJzYZAQKHH7YkEMvfXQyhYPNe96iWF6Z4/1SFaYfgSIaqrsi/hipdduJ7
E9GirMkQfsTdut9B3wgPqFLcFeSSl04bEJiexwDwuwBBxoYoMWrZP1o/C92f2J3fD+w+YDIIpTfl
pV10Om5SC1CU8c4dp56NMU6Aha+NhScsD43A3C8CYkwBDBKaEd4nRCqTcZ9iwON8OD2pxcKP/iEH
t84K5TuMu4F2DuyjJPQIsacMkz7zT8yswuSXwdZLAh9Rds+g8n6TT3dmEfHDl28XU+nu1PJdBs1l
R5WY6kuW/ZHAymKIfAz6Hiqx+ha7dW7RKu4oYt6cuo/ypf9TXFQldKBnMRnS30rjpW7s3jpzp01+
l+qKH88aKf/Uvg6+iBbf+/qgliZKgTdN867BCjFTBiilI88cUlL6PP8GXvMc73YMfBxmJdjkDAh5
bALY1/P4pXNBkr2waeztxDimahWSzJuTM4gno1P0+OTRzqo+di8/bDDfpHhXDELTd/SAlOmHjmkJ
IVpcFNl3QLFk/XzaoeH12GmxPwZnhvi1YgBlxnvqR0VGIDIp2COU2FzQlo9MSXbg8Y0x7uEQzM3s
ACC9O0vhD3G7LbICbWxy9cXVrJmZMYYPtGNkrXMVW2W0ybQMSvbNIsM+zptPlNmbUcCfHocsEypB
i2NqSPb9+gBxijC/4Rstd7Uc9Sl1ieVnU79Dlu7oj07fkXlJWz6Du6xtBFoJMU15lk8l5hBH4QnQ
HEOHZR5h6AHw8oWErwWTvCoDiMBxZhvTFjQjERdlOmDpbeRLEl7tIEUvci+ksvw6i33zbcDhgSUB
4M1zODMDrdKfR2PbY1LZ1pLcxywYK7v2Xb9hzD6djGnXG5ZMZkXp95TnnXg9LXKU3UEDAru/CPcy
CLnIkaogCknpYOMRy8Tj6l/cw0W8+m1MDYb5wJy9L71AkOjKn2gRRbfcwItlPpwamwruwAwNwTgW
cDe/gQqI/52XEGJ1EqngzO+hEysB1f0ddnr/rlhxXvMPST/VTirnvnlTcHtxwwlgjX7t1LR6r3nl
3POwOwrDPUBGViRnUUm0ZhFsCM9SHzm1KSVIHbFtopR180tr0O1k4G3aLOQuh1RZpbMXI3HDrb4a
EmgiEUDkmFOsHtuo2vaS+a8/81tgeYLQ1jk37GL9XuCFl542owIivP5kl+5g8rxwqK5e0XEHf8jB
tCKXZ+2AQPLAvnCyGW/NEhrzYWt9gdYaTzm3DHJ26AyO8fOCo/OACiUSVpXgaikw8fkh1adK/IMQ
zPySSEdByU7P5BfQaZgT+e5U8nuJ/4zo1xLjotEawSVeit30e8BeNe69hEHyGHudpoU/93oIkGWT
E708q4+cI+kaOxECogTEHO2LdxKE/ALc/5c2WY7WmLDsz8+gz4rl6OtEO17f5nSMqMO72EVrW1Mw
WhIJzAiSPFB1XtcsloyfeCmW3I9h2/CNPgsiKcgP91h/5WnpiGoSqeOTv2c1QqbuVtumojK2ns6q
094r50WvKUtTts1r3GrR9rSH1G/DEiJ3t/vH9u4782CgJI1+AuN91pOhXmF5hfjQ4kSY1SrsTy1/
MaNdjZKtkKM+rB1d1PWI0KTy9QxynVXBYEPBPOLl1J/D0VeefpAdbAq3bAuF2/R0AKkClQ9bkpBX
DZVnloxY2mO0Q3SGoe5WqO3KTQTkw36nsQKJtW03oVZHpJ6guB7Kj3UgUZFvGMelk+uZgFe3xQC2
gsCcWltVChz+ZbGnQJwAsWn8Diddb9NQQ7pFrmJaN6nnT98yrQczCFb4+c+8A5w+ldgImfGfAB+q
oywa6Y38sLkTPgPSg/GZAetm3+3wrCqe1zZKiND248jNjJvAeBhWmfC8/GWbc7KWJd3aRlO7REcn
5rjBSLyeAfD6BuQhGjfphT8EdsVyxm46WzVd9T+7LEM5tkaAyFELuq4wIs2ZYnhEKrK1xKraMVrE
qdrhbxtwzoM+eCD9EaQ8r8JcOTI1cZ3UmdBz/GFZaSVTVrEKToEE9hTMWd/9DKbMU73kXiSI1VhV
Rh2Jb9G1RoyiFdRGKNM7qNqX8bOs9oUWHEJy4K11aFIjDRKkg8RANSMkUEFmp+UrLo3vSzHZ/6it
EMVaI1bwJPb76YZswKD3PtLav0s9v+Sq8c9ev9QR634r07F+l80nAqwT6VwGx1pwTfvv+uHn3Q3s
m3hJOqjcccn2s5xIZzX/H4wbuvq4Tk9so/HcUdkJmXT7tVppl/kd46KgAvv+4F75Ezpqn4XA4nE1
IAfppulA7WfxtkM7hAe1LGuGLe+El72RQxoMQqiOFzu3HkzoZ5zejsNZBHD1T227XQozKI7vV22L
9PhtfeIXYVnbfTMqRNV/39BATFkMTz2ZypBGeu9PEq6JpC3ElgvfRl4l1a9evr1qPwEwsqil5/eX
IjuZGFDYID5mRl0Ko6WBmbHlde/MZZYt/aZjJXxwYqZEeONt3MfnOaPjzdC5UssHNsPb53pPZjFt
tSNCcMkZtNgFt4In8kn/t1YSH2h+qd/fjyAOybju/saeGRmtyPlE982vXFY8/gK9pt4u8nF3tYsu
An/3SKXVY6Y7vWwCvMmlv8fRHMv0+Wxqr2tYRaRfPaHHOwyEHJOU8t4T4M0pfNJ0uFpcTCXBzkY5
4YO4nRN1dITGNlCnmKMPxfSaQmaF4PzxkZSeRh5oPg4IDL+v8ZvZMBZ0mpuDxRwjVIKiposZ19Wj
6DWT4nRiwQzUBojkVZqy4QjVrEc0lO9Yd3dAa+09x9S+Esldvg+mtNY2Vrt/VYAiZHSgV5eohbh2
M/OLF4IAMyM7FmfninTG0w0DLR+t8taX8w2wHqDSZIgfX5GoYvm7YxPRQPwRZy5PsuQCWVW1GX5C
ZOuxuDHClpZpBteKPUPADktNvh7JMRHNQ1oSynjflMCQUaP+Q2tWCVVu9tyhTzVciyhuSZP1jHM7
OPXTsJj6idNSwnIhxyjgJpgJXk6ijnOSBxqAc49hJkqXpyTzqHT5S9vOTzkeU38gXvQQQofsR/06
oW30FVKY5ajtx4PxrXlBWEAQ7eYKbN//G96//448jAPegBOYjlh6xdYf+ojeKPY3eyKiupifP8T0
f+Qfn+Ep+19eDcj3DRMit0nXzD6CG8kzVwyow2QxsLZ5IGLtJBoq9ltgH7PfHzpoBO18/2AErxlS
Bo4Vi4ztTm8EOzVfZbTUhSdC72bAY5Cxam8bS5ppSiniQEr/cDvoKn3YYKSVOY9776omY2X55cJe
7+dUBYY6m0C0wkbLDOX8T1kV2BAOm7zCJqaf9wtZdbwnMDiMuM6qcBw7sTkTJM+dbZFK+axn3Bes
1zZJWUoYaQGksb3ZOttducSCShHqvW1WVwt1XjU07KgK68YxZ1nSKb1jkE+XkD2lehdQky7AWMIx
aVho1NtH7MGH3fc+7e6H6u5/sczJl6zIUGkWsyPoILkF/qIUk8gwy4lXOyGeXfrionLAfzB5CwpB
LL0KJJdgSE9cxBQ5G9H3ODXpNOJsAkX34ImyUQ4efPFlkCA7YEVv8ENsqUG0oKYRiZWG8DgoFF1a
uATmfxSsGTLXeY0bNUx+r+0/hnxPzo/g5c6rl8em1+45GZPzRTKKJ23k3PEO8XUynIf4JbIGfuiL
Xr5I2dcn05M+S9MKGiDzQOfI88ayYC5mFRs6Hu87ccjZuA+oHPn3tXNTakel9AIwbY1wklnIFQbc
5ALEBph3M2O5BNCNJsiQXep6KU63mOTFeyzHRmGBeDeB+O2Ga5DYu77v5KCBKXV/IkozWfgMJO0U
AMtZ5zB+4SzAL3AXoj8hJUInbnQmmfGVJCfrLHWFcW/iX3mri8EI+wz6FdpJ32+coSaYZFnqnhhd
SJmM/flscwTZnze9deXpo9JqCkCQTwRYwum5KCHZ7WubaxnhtI1MhEXAqKduTjPLJYMy3JBZKy9r
Vp6e9PaYgZ4aLv5fWDbYWvM6KoXh3wQb1eKCPb8GdYLJl5bewF8yoZx7zc6/LiX9wJmID2aV0NiC
cflwzIT5Ny2mu6tyKoQjD6FI61F6XapbLFVMzKsAl73xWDCIDc0kIdtjCoMU0JiqpqGYYqHmrS6t
8yeUKyFUQFvWLjvu4VJj9X9hp/1NIi8EcrrZzpB1On8RT28gt0b7VPBcNOPf1VfW/MJ7JYiu3aec
zJ8FphqoGIAnDG6gK51QrXzBh9u0Hdu4L1wvPKum00Zq+nCzFblHU+jZKFzAu029o2LTSC7KmWLe
XOW+C9U+j/Z0uDw3EExiz23Bqs8l3GNVpVf65PhA4WFuG61N78kf2ZAZELsZu2o719liXQiQ0h9F
6sa50aJXG0t/YqtRuOgtfyQYVeN4j8DO0oIoKhKKBztQqFbPxj3qEzk9HHiNOgn1OSIwL+Aayqos
CXHCbSzJVZFYsZk/OrbftoSdYVXLz34p0cEt4ZgnONC8HMwGlHrAkjR7no22nlxyHhe2OFG2nHZx
mjqUo6OGv/9C3zzERj8wzObwY9Cs88MhcQQWPzkSKurHI0gqp18gu0qoZBE+irORIkG7rHNz7jYR
8oZEp2ic3yrrX/jm3VIPbFuPDUm9SBfdTTs2LhES4uI+yv4AcSs4kwTpIl7z8p+NuOdm7LQCG2wT
R+qFieAZbiJMmpyP2uNGIg8mCv9hDF2KZ+R8HrwE/HpmLeahqcYtk75GSqdrDM9R1TFMYJlKWfux
0RzLp++mVWoh+pbFPC1mUe9r/BlVci4sG57bN9pB1fhaZ/QjIYJ35+WZ7sC0w/jPe2ameneBQEef
Ic9N7YYU03AAN0gDmiN87Y+zsRXZXbrXaUHgo4f8usv619WvwSI9Y2TZiV5FtJcMBsqBvme7NLBC
pIFwdYAAWeDb3Wr8eZ5+IUt3EP6vHHEaP2KeqYtsz1yXLS+eIQmY1ndlEWXYr0mQoxeRNAJsdFYg
g+VE7RZxIjeJAiIdNrG3md/9ZYFfawSjaKyUhiO32Ab6for4voKsRfNLhkDUIv2Mf0tnr5340NgQ
t7WxMNaKdUm2tDkgZ6Fa/P3Nt04mGE3/EZQPRSkXLVJ3Sm7BTqe5HwGGukW4I2keur+c8FRiJE0h
FInUdyCxPuKisQ0zt9xuLVC+OvIAkXE9HwM+RzaZoO5FbRB78nANiDVRv6E1GVTkFBkyf9dYv8ur
LeXODX4pXVwF9XK1FtrUkhd2NA+j/wbb8b4+JkOBMmIfA/WT7jHAFNJaP7QA9aw8LVkSqp3gZsME
PfwM4pe48zcLoNT37GX3+qLMFnvyUeBhiSCdCL0MPAwhG5hekyGJYkSSA+B8D+IBK45w7jIxVB5L
XL1JwC5sOBsbLENRTcTTjGFMwPl5taE0UKweevwm214SoPK3n0cY26yfkFnYlzKpMTH6ayyLfg3d
E+wDCC5BUEdMJhfdsiCjBD+y7AgiZaICV0OsZRMm4cXfRXyQiFUFsqCEfTEMYRT460djWHuNTCg3
5wOqs/6s6bvdtW99ktxpeyVdbomIRmO07N/i/l3MIJGuca1fspAe7hY6EsRfMQVTFhsZCA42yZVl
wYclDIHe0dV7co44ZVpTkGME/xeyHEtezmsGkQ6tdfOaEgsgD16kLbjN8x/VqsQwjPDx2OFOZ+dR
LUvtAfHva9a/5fhb/wiJF5BGQ0FVK67p8L7S1fNih0sC+yT2bVWBX6jofLcP+qmmPI815kRfPapK
XPjEgOJPsuJVAiDU/6vOo5UD/9yAnK00aLvr3ZgBxBEraL5lE8NOmz6X9m+sgKaGzj57aSu0jEJW
aiINqpBfvZ2DPPk0AWGAOo/X3YJZjJ6O09RuKluv28u4HzrzaszElfOjSd3vshbbpumDkLIjjBRx
IPn0S7SJNY2OWq6YkLPhjihJLvscMOoCkdagGbLQYhHRedImXP7kmi4grHhl+DgNRTRrH/GrORle
xy2WcJZwo0NE77FbBemm5qnNXFrqMMmoWslgHYVN1U0DbxlPlhFDuN4J8DQYxZe+qBHlY24lFpfG
CIi85LahR73eJz4gHr8gVxgvX8k/YDCRs1i/RdjcCRiZg4QIG61V8UBC4OYVc7f1uIgIRYsPpPZm
1kojOHnbiQxmoL33iI4P8GRYomR9z2H/EhsmdKHvcn/9hqdF8gxYL6wQosNonugeMKRUDRZadaYU
XNS13rvPZ3Awi7D+lSwJbNKSQdpMk+AU/1ZK86k17gGrud0oKywutxPqTB+Z7S6XkHEUC7n0EoZf
j64pFl4wqShwJgZNOxIiH2hWmQ8QVG2Fb4T/P0bpClUokUgVcDU3ih0wGwZyYAF7u3gNaMwwP+y9
+rOk4wfEWaNTA9UQQWBmqJPXZUxPJFxct2C98v+V3+anzAX3Bj5ORMszOIN+usAf5vXiCMj6fl6D
CD6cSNggu7y7kSNhJq4PGPDaCX0h9L9v7x9mcZ9yum6RxfhjvP14GhiDGGHYPdCTLk8ZW8j6mEut
cfpAKvB9tkWAjpPgIgiZXoKjcoR+He4XNGlg62pzgc+vfh6YxbkZAnWQfHeMZ6d5n5VCtpc8sqgl
/SjLhOyI93ivHtpbHCK1xUgZbonxwiQQ9JxnmhEaAtwal8p/6FlbopIXozFrJTu7TiZ9LL+46mwp
tp0fNrLaQPjSwwEJhX6w/4+LkoaIJpEr03ZDnqpDcRM7zj7XMcbK6OSsBu3PZecAnUAzVJR0IMSt
ZjvKhr31dvADIZT1VJkjMLAnIpN8w9N6TEWzLpX7B1qsx5FFRylBGjujznC4b/D6h0/n1p03Y/bX
cmUf/3CBgSnLsyX9YOofHcXxO/Tv5HLJMNFk3gwoGR3nmokk/6vdfWCJe/R2UiU5j9KRtc5d2TLa
i8egNDy5bCVM5BQUgjjGgibe6zfo/ntzuiLyFz4Bd3Y3wJXvAmWPIBaXoRiiOP0UmcaYiP/fM/U7
JJW+uepSE6rfP//XGI8kv4+RHApn/TzrQNXRthMscaUzTfAHvKONuv3VhXHZV21Xkadx8NwABN1v
nvsf9uYAj56p0Eb5vdtcP7OWnvL8z4vEEx2DIEGzTneklFbww7cb5GuM07bmkD8ViX/Khij1474P
8OuQucnS/5VYF0Ha25Jx3doxoFiOINGpNW0KSOhwzWGOGN5WpYpe9umYbd0937E2pEfQA2NQnPjl
TKRHeJGbggQJFEaFAhLIqGDgi4p2bgtPk4UoYt0Ah8jNfmsyEcF3jaTtSEbgq3T4Yt/8i/oTYsRV
pghuOoqQkdOjX0FSlf0riEObRvgdSYWC6cJ/miDvbm73uRxcW1jL+CbRWXyybnTqK0fjDDk1TOpx
dVf+gobc3WdVNt22SlsehEyKdVCmaAp4Y0e9QX/0T1WFzybMqUVeXMrIdvWCCilsYxWsu0wRLh1l
/cn4CsdNsBFDq/e1QS5ssfe6WPZ0LzLpvlnnSkfJW7NniKwtkklJ0/RrSqJ62KWpHyesiOGEg+78
+9cH0htQ25/u5v31wjFjS/IC/4hC8l3iInIkH56lbafoN8ghHVBnbX1tesFq8Vv6eedDxmsV+4BJ
LG6LN9sv8Xd7C9Izky95uSTfathyc+gpVQ4R128uNCiinm5DfKCwfS94+AA62lE+CGWQTjR/9rSh
EnjgTzNe4bgaGZBl0+nrQ9v4NeeMBcnQPtMARSrGIGh7svQdYZy/4rd3bMwzp41OHgXaWN61LlKC
+DW9UJ1U+U3hb7AyWFNAXTyNggxrW7hLNR1DgW3Q0k0Hs5b1E8ENxq3pqgAjHwWPtynf3JOu8j3N
mndBhbHkEGc0XuGHGnbmzMpfUxQ3GzelJetfXZldNrs16GZFXUmQ7bpXVnQM6wBezVNZaCxiL2zh
xxAj6JP9N//TV2z8Vtqdg4ZuqoFIi+VoyN11owhTToEs4/rmd6VmhKNAsi4gXl/zFwtMwqRpdGBj
iK2e97LywqZblFdAD+msSSWHKv3FsNPLOhQuOhTzhYQAy7lgBGEhrLXozmsuJ+bMpMCBRNT4Qk8V
uj6tf4bdA+hZZ26jR5IWNwdmFZmPy1ZGv6mHBRY3v6HeSJ+8qD9xydFD3OE2sElaIv4WHihO3hn/
4hfb8Dt0SoJsZ2uDrKOoq2xPX/C8B/FWwszW6xX/pPg7ks7FIA8+DrY8DJmGzgrPcXpEKKnr+wCN
LZlSOuA/IR+ykYBLV5PoRBARUbdh/UBi8wTsAm4D7BZy1m+KZjYA7OpQklF46FPmYDqrWf+0CiGe
qtbYkfiNneGFc47jBMUUJMa05Oz3cjygTPmpXhkVyRv3/FfnnMgANmvQm9Lj+JJBjFbGGqodxCmJ
AFVVgLeAT7O0wsCyDW2irCOsglzS2Mh0kffTOulHgUI3/pQZ0zksy9oKESGUpBs82tpjCz8LQjVZ
4TB96i0+GEaDWRZwj3U7HWuJS+5ll16QPF70m2oWZlMM0aaSrkWGTG+nndHF6X3FWs29YMOYdgLB
OkRY8WFhbUgM8CBCNfEN7gt+qq+i6ZifuFAvvZ03TXe9AyOlmq7uzyd1/dCDhacv39pYDmJVeoHn
C9D0VMcXgWXYNbChvdqXePuUmkcpFkBKXH7tTMoyKHwUZIK8vkpt0nRHQ23rDGjBxDMQ3JXM7E3/
dmmnyz6b74cUTHrNWme051d/2FkT6npWJoN+z5ivvPX/a5hcfBeRhJ5IaD3UiMO9Yyx3W7oyMUPE
x0oo195zrHyt5LkHwmpbC/NORFgtH4EbOCsFBXV2QScQquzQPNHamSmd8tOqw3xepouNx97GgFuo
eSnsta66ynt+Mb52sKpGOEriqDsluSFdXLS/Q5y1qTPe+/+mrHXOc3MH5J3JNet9bbsCIXLT9/DI
6ewRReHVBK8NRuPM7ca9ciMc71XWHLiOb4+h2GLjTJCBadyBq72BY9JlqY2YKmnayL2VBCP2gofp
HfaExdAdzMhm5Z364cH2XNKMlYtsLOYqpTeV2zO3NVeKMvBTQr0/R9idOnlxf1ZOs/dkQtWgtpFj
E3PIGlDeTbzRBcWqWNp7BbsvMVV8bfAur3grVgSW4rYOxgjkFD40+siTbL6kfBWUHlrKJWzuTcu0
1K/euQF2AGXYBSkn/WX0ExUw/DlTtB5tuC6Cv0gFiPSseVKniXs+OpTwNKRFMrTHEgE6P85uB84c
4K6qTwRf3kXKemJQrmSh2RvmfbPvQi4Z/rRyJy2UWeS9AZUa+cL8tD//r5wFJG5h9YMQB2hCb98b
ldYcxGI9IVR/gNxPZM4We3VuuycWuJmxwgsVqbMI9KAD67ZvhRkIC5UgR6QD35YI4yVFEyRmCVKr
IA66HCqKY4eCP4K10/AlWIxl97qNKxliRWBIEkuqYu7UTNwIKCzTOnLy2RSaMFMoInap5xmeaOTl
FBoH0Q8JY4EQ+KpQstB7lNbpIZI5+uHNtK6WulkByq6A1E8M/z2VvlsDzzvU6rb8Kh3K56hsj4+1
mIKK9mK0/tiq6G/qegMJLtpXNKoICH66htB3S2RNRPym7fb5scyhjAP9GFRwRjyHg7B3PhMbnSWS
+hPoxjhrgInn4NIiFPNq5+HMP7YdemaF15EWs1NRUWoPZkIAos9WaGXZSyHClxxv+0SqonpRL0rU
M+jAidtgIgHsvFLF/8IRfbpfcVHY3nFNwxB/mlevQ0KNbO00p1ckBkAvX/wALo+/H25BVouNIY20
1bMmqzGodQy2mwkR7xwRhbNWNlWWNuEUOON+BEmp/QHu96jRX1ikU/QgWfKYmzxyDOmmzdSIOo42
blYDrn9khCCOysDxRsoHmH6r6QJgfXFPtNQnKL14fzVO1+pzOIn0q7LIXsBakHyfWhHCssLQu3r4
gaHrqkLoWxFYd2rWIfwkvyozW4QrbTUFQj2JYn3MiWSBYB8q4TIYWmx2CXw/jJGbDoi5dAZ6W2GZ
Wh1KQouDzCSzoDZ8enqY8x8TK60tpGmeCxthDi8qnmrxR12E95F0UurNKdYDKnwIpYFXZrsocjTK
dMk3RGMl/KUId0+gt8ZqNTj9D1NwdW5+Hnz8xkWXGTOw67vuFv1XrY+qUPWQ2gK7bFRAo8UkkR8q
Q0JonvCKK80LtXMOfgpD17we0QFmi7Zmwn/R6Oe8rhD6rn6gXTso8P1CEUCCjdwgOgVMX38c4ZAV
3dI58nbWO/MkJPuHrKnv6AhdXbxQqsMO3Rr0JFGq5YeiV5cQAIrxZdyDRsGe/MpDWwQC5K3fusDB
BXYx7aAKzpG2CvcjXs1z/nqyxDjBn2Q50nETE01/EWFQgBS/WL+WR2LgykKLMU4w7Nj20gS3nEcE
sE3SFwuheDLa3djsVLijBqugkeOTZ6Q7YqbbXnqEdNe/jbEqUHpYHz6aZybKC2kFm5dG2sOglQHJ
e0iYAvrT7sXPmwLuXuCGezr1xKCb0PkY7Xohd+wG1Y23WGHyW/8mDlvRmNVY4smFLGbGF/xj/1By
W69G4r+Kz8uYclZsIYdbnZaHIMmM4f/jpZUL87+lhrnO45n8LdMrJvPhDpTuYNka20LbfXOqJxns
KipyAMy3K8d0WxQQAanqMz2wU04muD/XhEYxPoHLIy7AtSHeRXB/Vx5sYUndHOVFuNLO6lVMrFiT
oPKZsBi55FHd5+fC4lL3eNHtRf8q1/Pfxs8HZ+hysulWtNk1A5mgaNGKFUkQaXM+XU0UFZv3hJBQ
HM+0D79DloCtfgkf3t5/RBlGtJfsPsTgslfTBplGBVifEfgVxbvQmCDQRicm7z7hXH3AXfiyb2le
e10LoYLPKjOyHsyDbUPCLxydalNkf1xhxRqD4Yog6wU8cVUPSJiEqZvhAbyJQDGb+cCn0ubzd80B
VbwYMNLzZqzRoHtSUW66MBlSxwZq5Ddd+oD7HkXNUUma0/2TXFZqRXMYfGGzb5yUTaf7iCcVbCQS
qAsO9BdhrPXgQqDT5/QWXcTAUj+8TRb3ElepVTi66HiCS+atAOERsiYhrMFQF1btyTqudHWMKRGF
M6DmjdSh6YVSYE5qfrLwxfNr30l6I0txQ1va18g+cIxpFy8sr5pBo1HkJyIiiwE2AUk6hWkGE7xc
vNn4xeouvEqowk3l1DbqbrH5jJVB+d+Zb95PizQagno96W3s6St9Hkqytm93hAmrsdMgPDXNveUo
+iI2vEwIF4sU8Hd7aUrp16VJl9m7yT5pqtOVEOJCxcIsBWGJMdsBhwj/Jp8iarcb+L+EVi49GYsX
NK8H643wx/C1KrewE7NjBWjbBSzmsjVpjzCLFmYv536igUO0mPLCaOdtL9BDoPbSDevoRQE2w6LP
mM9vk9CuT86WAPYJ7VU5KtvIDeo0ahIQsmAvYsqawaPhmHmpXYjifmEdxK+ZJ2f3dYV5Br8UFDwQ
pGYctFDb07gSTHrYnUaYnQMwLpkPHvT0Rn1md6lRAwN3KQoWoFolgCYxVKa49cBIz2/QnR58b9K2
p0AgMsiIqu3hthQmV3tV7Km96abY4ufmBB2Vk4D4OXIxTsGg+smGMN1jRy/Yh6YGW4GbxHD5FRTB
soRVdIEtFSkLQW6uH2VnmguGoLjVKVNwTVSi/mm42jWOQps5J3QQhPQcCyAlYv/VqF/4Gc5dpdqm
yiB8jp1Jv7nx15PyTsWZDE70a58tgaIz2EqMCPu5XUruRxRj1B62K9l5AS4e0LgS7xioAkwO62XC
gRrNJal7KPiF5pZTl8u1GWaq4hxkbYPFeUnVpZOx4ZBTJgzGPl3RDrghJjdiHR+KeQr2PKi2PJdy
mpCGGXImBSkA6SpnCrsAdzgvDNhBEqLxKMqGv7N3bJlcKHRlQYgDMm8tBef2FdHLXB+mWkVgPoqp
Gb8N6+B5Bn9YRV4okhmVM9c2dEyPcTvaS3IAHq0tTbjZGcr6jPTnDUntITaKtvvIS920ooQdtAfX
GLgB9Quorxhm5oxXIJDOXC2G5vxtG8IA+PyS5+vPe8HRqORCZ+HxfVvmB/r9vkvBmHe2duOSjPoX
fbL9rSfi6cXriAfWtz7hRBLUT3KvvualAKgmLO6Ul5ebxXoLYmJo8Anh6pVrqz8W28w1IX8EMWZh
ejtXqaMSwbU5pLDWETql6D0cGKPICuJU4ii0su9FTpZ/5bcvZpbCnYNxJm43L+ttwWKNCozwqT23
dwAHDVGiBSPccfa/VaAmh3Lsids3Hp6IRHpE5n9NR4D6yOVyZlyXpmgQAQDfbgTmJsz561/UO5/u
QbFmgBndkEWEZXdO45WFYpGqnThnfTcyZXyMEgl8nps5a6hqa5Y5nciQH1W3/zh3ka5aWf4/4+gk
qEspQazlncc4obnDNIUJQzLbFzBNLP6rlEwJ7U37r5zb41ZUFggdPZnMAwSZn54ARh/9oqBn9CsP
ra/bAizTEK4dQT6++peCUMUzcq+OaMrd8kuyFIFjvG5TAHbHWvKzzHPI8Wz0ch4lq2x2pdb6SrdO
ykVoNkXtpblvPzpcm9OVHZJqu00VVBRmV9IqFuoNWDdsyYmn4qDUY/UX7UfOtjR2ZdueCVjJnBB1
dC9clZfFNs8d/rBCBcBnGZjrbl8rxRImmbLgz2wrr1sKWkjfPi1D7RSFxF7kV02RDoGpe/R2A+La
tgFRcw5fQTPCLsKuc04J2IpShh0N9wen5GWxL81Bsl2hNQQfU3t7jPapaRZl2v3avGdA5GxhKX+v
Vg87nxytcubE+6K7/53r0BF2CZgkkXe6e6+VHlxrvyiJP+pUwtInJRvOKH8VF8KyB8UHAyzbTjb9
ROiHYAK0TS02DX/2dS+9/V3OM7FMZVrfVfTAvYgMyqScAqGfbrAGAMuMguZ9YKTx/mfouvy42qv/
xO+v11K+Hp9I/Brv/jKVLCKK2CEk+U+Y/eb3MDER5eOlli1IoV99E7D1U6T1gkiluH43s6+oOXGP
/4xJN96648/fFRxBUYCDOv78vYBJZA9kQCf8zFsrSudzkjjakHXSgDHwSRiJriQo3HiESeeFgCgP
xg3fGcCxuCkIl64/Ow9cj2jl+xMVkMyxX8FqLU2OP0ZSsA8+b/MY6rMBKuPgpsaCJeKmDwGEHJqr
d2ZUUctFKODDp+UnNWNweS0el9ou82CISW8o/xHD3VNeYlxJMeWIfV6oIBQkHB/btsFeSP58RLaH
eJoTwWtupP9GwOkMF6+D6P4EMUiHtQ6cwNk8bnPFfG6RT3ytrUoLETlTH23LzZ7ginS3uLGRdkiO
QcuXKP9gfFed8RynTOWezFvBL0ragzmlIH5TZMw9vCmJNlj7TzPDQZQaPCKG8AkCN4e7dsHbZr4P
J2Ugleh+whh7YGKXbFkUTQlDpkL+2RTetLmsr1OXz9GulZY74QDORnQOB+1MeugE0pHll7WPKFIX
8ZwJJilz+g/e7zqjyR4XqBTkvR6VHmERy7W+TgwcIihguObO52/2LTpSQfUfJkUlQxYg1oy2QCbr
lv0S3TjyWwsdZiuvccKiZT3hkjDW2JFkV6/AXnicUqC9U9kKnFkrT4VcPmvDgyM1Ze3IiLTut9eN
dSi5Ih0Hg6e+ssaeGTAY7TwEx+CyqxIhWFBOknI49xKglXRB5l5X9xsjFh3ZmUmMqT9NGdMmwZH6
S7SS22Gyo2u76mekR5eAmK3IZwJCmcgtwojbmjSa0H3pNOd2+AKQV5We9GHReABKOaJRrWCLEDN2
75XIWZWhVwhbkuvZ6h2H0mUPRXqJ3qYaF0YFTv5GQ01MzgDzzKgWStT1heVf64pT0F50v5j6rGQT
tdLPxqDf0xU/jD3boSv3vpXTyzLT6+tVumACPnPD8gkMy8TFsnkALoQoASQkFE7fQUCQGDsu0UTL
38EcaYR+TlOyAu1gCUQj/6+sWkwree+oElA55B12bTASNN+JtirRcwLrfBFke1Bk+oeH4w90Ovzi
yjOnD0RYeCEbfPP/R5BMtgQVDlZ7HVPUHjFjx6nx8vT02+dY+jX9kZ0boxnIICGXZGRvswfvDAMg
SMqIeE2bW3IMiOq2+EQ4dCn7O1kcfjNTUSRng+uOEfyXP89WYMFcOsMpDhAyPadcx/LS45pYwsVJ
M/X9ZixDCDTOcH+JSD8TTrpECoQhWwKh+h3Sq7+6XefvuPFZ+HLBlxssJRvvmBmTW1jZPkqj5we3
9Qyl/S1I6FE0xCcjFC40ZszT9FyuOXdyxb2xNymV0ILEd5G/Cb+avRmZd0rBYLCWhwiUWGkSVFSw
USoJ5A8DsW1UcfiXoVGmKyqUQpIAsgOUmNAbna880pWvIb5e3URFPI86OMdpdW5aYAEGks2JBAxz
MMOYtQhX9tu5cp8PiauxxXpwpYmow1IfjVDmxfhwdjcKd9vNK/qve0HyujaUz12EDyYLrQMjLOCv
4PEvEigggrTPqmKU03gm8cGUe2f2FJs/R0l9MULOB4N35IK5Zur10m9JxqtgRS99WxQofPBXEZLJ
XYmedfwtAVNiW9URX4MSJFVv4HMyCDqO2aFRPMO1is8hkVjegBHfwADJ17xv8b4uAM9LjzX0+pIj
+VfO2qp3V5Koym/aFqi6MJebHIhwG93SfK18qzRVRiAhHm8qgPllg1kcwM59c/nuVUOyrliwcpn6
EGk+Ig+fI1LqFjuOC3Pq900vm9uZbDjltHTrlvvW78exfsQhz2386WQenIDsfQiG0AK1UAr603J/
WHGP2CO+rJZFbEF39cxMmd5wmR72gJyGNyyNWf5myjxVOlhKKafLlPkGIDWNTcp3SsS/DgkjxkQH
qVrLdLwMVUkXOkgc0/62v8b0BE7KBv50JBmR+pJYzL+GjnFS1mlOD6qh1A4Mhp4nrrCwSkNgVO+D
9CZA4sgcWynIgobbg+HTB557oTGIY7js7BsjA8qsTX8vnnACmDLeQblIPAmNNlM6fCK903XctPXF
AUfrk7CHP79VBmQMmfosO+utEPetbaBlTo91Q5WXEtEQvnhjqDzMQd3ACYvEM2Yj5WRUX9Ll3D+E
4R2Msawaq6yDLEnklFwePJU8I1Cnu7Ga9kaTVL8fQtrefqc9mq34XHrv7D7n/cWpaDOKx83wEVgF
CIpVxiLqr0VMAqyXmn03CWG7pIEJnEC7Il9WUvUKDfYQsJkri3bQ7qzNhG2mJGjUa4MJlC7eccEN
mPYhPXls36bC3tzIcJd76TvDDs661kW+62r8pY/nwcl8E/8iDWi2WoPiyYVeDV93vgtJyhTAiVMM
XGUv4qnX8QlvNiALhx2tS1irikDIpixkRCtSD0BGW3AQ3iiRsSXOtkXLgqHT72y2pNdOe83EOp76
a5NbkvsXk5dVp2kgPVhsO3sJktELsFW0/pWUeEqfi2LsACiszH0bDhZWBboWhmjvICMCwbgO7Ncz
j5P0nuHmA2AOv/Z5uVOgUqvGv9B28p/wGFW1sjHXmept9pzFdfhqsddKFR3yrL1OFPh27wnQr3cS
VdatHM6if8O75lZ1je3Nkyrt5jptkOuS6PEw/UX8/zaXI1PJB8d9uvh42qn6EcIvPC0LrtEANEbT
zu7kzkheW9/d8f86VUzZdcWJKmD5efJSJ24RSJ3Bb08iObXbEK9RMELly1E8+dQRQ3NyQpubl3Ce
Dmo5LbtaSob7t+rW1G/b5oqfA/LP0iRdpIF5dfa+0/0RsJhb2Edg5axetWIXMLof16eX/2LXbjSd
2ziip/PaspGFUAluwxurtUQhbLYPi7xhYiER8VCMxiVAIi5MlpKexBvQ7KqAKFer4VxTxmEpZyfN
1dMFuMWINC/QPa1Q1+2OSPPAz98aIxdUnze2bLMHIbkNRVa1dClsN5TqlBi+yDOqVQTcFcSJmwMw
UZoHGBnLf4iKHbu3iLktlv/yVkRLf3tx4TAReOg4AO+b0ryGqZXZq2GR8/jhOmFGShwbLvhD3eyk
2Rw0D4YPnhlOhlmebjUywLohDwskwNQ+IEwW6rcBm5gzhd9DcQV5JAtfzNeZwVK/BDR1bkD8b47u
crABUf28EMDcOchxodF+kPPeEOTtYDfAAwBVRhp9vcPcLQn4RNxQXAXp4p47kSMpGxHHHkZYIMJ1
dcStVvTHzsXIitr2swMVlwyiy/q82Ve6tq4I+XI6PrUlq2jsJKEY0QakhQ2j3AnCpRR4dTSkNrtn
HcTSZJ23YXPjbiVPdDGXsbsQ9+KZ8B05BGN/o3nLwESqKSKwANaK7ng2ncJdLoIq9///KkuanKhM
XUF+5IorrHE2GN4Ial9HET+5RDCoKXlIS5/R0KnZ1xR4IzjNW30TKDPtYTlYdadqphePMvs+a85U
AeTLXVOxTjklUAo6GXMDfmJkRQjqvti/5+Yb8dJWTNDTLA51OidRSoNMY5nzTo3AerUkef6wU555
Z6Dp6Lt/R/KvFgY197Bj+I9Fa+S+gs8DxKvWpkY/2aycqTTcEcjIcHRcGVRSWebuAQdjQPJBTO0J
gyDAYNwxFhGAZaS7ZTB6cEgBRJo9E3GtZWGLa0bLypbz4YnTRSFEbWvT3unYtnPIF0RXiu3iHNcQ
Ytfz+MBe0d2kP2M+LR8zmOaaGwlGAtMmbbzZXAXDf8jYnCZulElBbZpbbqB/DHek4oS5wOIc4ADB
vcJI3boTcCFFuFka0rfvdg8xSqjOrYqGqKnDw8U4DQCfZgy/MO+zixRhLDelx3LKXr3vkmv48zTf
28TAd6pqcA1a32PBqM2VoeS6IzrUi3lfdeqyyEiNowIpcQWCQLP5+A3Rcjb72lycd9t40quIYy7p
DJS89u3QUIyIX2TmOoLysKRsLr/GBaIhJ77Hq17ibk6SHX8SearlRZ5gOxJzmtZHpoMDdg9V4M/V
8QyP9sv67aXodgBfjA0GPYynK2TtEDsktmqh9u+uugJ28bGbVRlcTkQuVVCpRvBU3PU4G4BFeRTX
L7uPvDM3KXzRMwwg6odRXTBFKMfhW6pOXUKlKSryBvIBtK+dwBpZp+hkxeu6coidX3W1i1pT8ee+
TUOSeot7Bqg8uACpLAy0ylnkO5io+Oky6mlXuEtXWcD7IUBnCpOD8BIoVOM+BILy+N++9ISEENZ+
aA+wsxEZwWTFC19BPyxh+xE65g8wnFT2OcS99BcFcCTR8Mv0CuIXMzLo7jj9hZsdxjG9SD7tZrB3
I/ud84aNJuaQRsPfXuEEAdo49U9CF8SxE5ykMfcyjxQs5m76efHRO6qlTGI2z2oaPCXyUZ7Wu684
sEdXYCn677eoepPtF8HgQyBJ1/pv/5eZh0sYqA4rZsk/5bx8z+pJ0aMjrbUjoFERwXI2TyJuEdHn
AtbOpepHEGIvSu5nyhG1HHiOvKB95tnNFZUc4jx+QIS2Ci/NTfeKSCZGJM+zifet0TcsEGC8DodS
sKeT7fJh8v+TEWdNPPXkRlhje5cAQVNztmP1mEdSp3GB7j6M77aUggSVkH16qxnGTbklDpQcE939
Y/pUA8M+8wq1Jb+OBaOOfaAtS9U/axMEZBCF21ijZ3bdkHyuEWqBvjqcw6SVH11u5x0HZLwuHf8R
R+vzpIgyGXb1TsQRaKY9Wk6AhN8C+P/gBAHsT6GZlNrDcz/3cXlMkhN4alwmcuOBkXf09/sLLtWO
rcugibDY8G22tBv7b5OWJdylT+OKqgROE9cHKlA2e9YHOonZEaAXIlvXsqpc3smQ75VD08HVO/80
MecyNbr2gUz8qdE6hVyA8GpBKJV+s9EC7ZYIaC3dDOH0RDJlHxmiPlRy2ySmv1kpHCxZoyGG0NhD
B94p4AQpOseLnQ+6GLpBm54k3hhXwtMkF9rQTJPbn9oU7L0OgTjDO/yC2H6ksSlkNkHCPk0Rg+SJ
yaLhI0fWCsTLTS45nz5GyRzY07IFp2o6A68GUcPryz/9U9wM1moWrqQnE1JJDoK9yPpv/cz4eAqu
4gEYZ3XZeN1pzm9SfyHEm0/cAHiR/djQpQAZ0A6uR+aHsMMqd0wtFh1YhtruWGitU9gablMxCI0c
GGepWP74myg0g4D4LIHF2TBTIq8ha1LuLp/zDDQwnEsvdt58kOUiJyrpXmTTBVORYkomMCR9evn7
1u7UI1kZ7P75Wm5Erdd3w+GZ0mgMaxvjGe4xOhYr/C2q26sgFxRAXplgtrlxcZyLHrM4RrGhzD6j
DXnyh8PJ/z5WJOoG6ORikMdvO7D9w3spg5zUXrjXxwr55k52DeAGx1wzizP/V7TLpTZHpG+sB74r
M090kXoWa8krGDybVficXHrgzTFUWlMEM4OM5c/dXZX3uE9FfYruv/TisJqlsaBaRl/3geNr/MU0
qBOyCSIt48oILxzMYa8FrQUFi44mKK3t0CzNZNdmjl/qhmu+tVAuDvZ/9/KM0hSWdpVXiptnov0H
ifF8NZ9GZAZpTOhcqOTgzcZXa1qpjzNFzRnwMWWcouQ8M3cY1TkhoXOE3VbPYrvuAM0nXF0P7zZf
3o77AayWZvrj4511+FBydXHMHOscg7kkvzOS/q3BvfK/nds0/ccXaBBCwVJTAcekGCAnXZ7dTMss
ebQF0kvALNB7hZYLf+Meir9ghecSmyDQ4yHqygNxomMunIJw00mRxBUM2hoz1vBh8EJzW/k9Cm8n
0L9cZ/BIl9WZh5lhjmREc9diD2bSbiGfpGsCAFmQrS1tkAAVV5j9S1WvphH6ylqQVjYm0tSgRWbu
wsV4sUxExy4BCRRuiqhAg9GPnYilK71ZUZEhjbSQKaSUFminRIYbvhLE/90wACgUiToHMIIg3jN1
xOX9di6qBoapC0SGglCMbxmVOSfinQKDc5KCkKaJAyKMkuyTFs01oo95Lq0+KenXQTzOiLwyKzDd
tqnAQWRVyROWFt69ortkiupqfA72d0TNnvMWz/Tc0MBlkpRReezKbi3TGnXmUmiOalPejhsuZxCK
W3suRawh+WxxfFesxhWp/fImhFmjnLem8TwpBJpWft5mxsNYh6078dK1LpzMu6k3kqrAV2fOAcML
vO/4F4Wm9TdRf41JFFEXnR5kmmZvVn7Fd3mQQq27ExRrbQGTw6I5qBwpje+56NyAOPRn58249NDX
/FfyoCdeADz3wMXfDv0NplSe+mBkAGz9huaVGhSuiU0kKWOw1pExwz79E8bTEMYjiwZrOWaA3p8p
mVep+OJZblXo8DSqP/x9azVjO0YUuHJ2hmQ5/7b/FpE4AbgWsBbfN2fbS2D3xaClRVk6qHWaxElQ
Xf+FdZ8J+YXBhn++6S9n4x+cyM5qyAjw/ZJ3n44NMu6dbFV5zOKJIrP4syapv7PPmonEK3/6KHg+
MEZXYlXXm3TfS5eBSCFVRs0DAkqI2TKgj/Jkg0zUb5KwggyqaFFWfEFXBv5hniPpm5YnGcVuE8xL
miJ10l9m5O73RfqU532XEcQWxbyWxMO50S2ChF8VDs/nAqXce8ZpXCLtFJgaeHXsRHVjdl9J2h9U
ctZUfuKfRCjTVDIqOR/1fP7h8xFaLYAUHWL5IQVvwvOTrUCtJiG7gQUFPMOMSerHeTTLYP2OrI7n
C0SZEcJxd/fGUL6+SQNRcMaz3bcm8uYPBN35EMRKJYumiXl4AwVYUX1CKBLb1iWtBvNQhJ8vJPF1
YyKasLwAzruE2po5nmpV7csdA0h7rfeGMewQYOJG/IsyFj4qqEcg5QvhE1aNkfmg1BsMo6AaeyW7
YPDyCzFmjYIueJREJlTvXWuP5R06F/PGnkvnB+ZOUN2js7ompCT5rZ3BlMRV+QSeKOxzuU8jPpii
WLfkJJMEK/LnlbRbPa6qfZFdGb3jEb8QCH64Vj4N/uHsu6+JOtOU8Gb7IAPStVvrBb402DJEfUzj
NEl7UqxT+Dgso1Bamgnvc7GonYao0KYp0tZlFafOdRyxOKR6Dw86SaBQSKSCl5CMZ21mTEjt2pZq
SDMyVkzI6Qwiavbd/8xLp87+WFQw8TkGTf6J2O/30XMiuPZz1Deg4hjmpJeVZDXzuK5Lvi1VZOQO
GFEqkYLNpo4EMCK+aK7IjTcvzzFx1TBGdBZBdjFxz9I1Ty9zHCUOLn9hFYRRKM9JdRCN+Ee9mLns
+ySs/aqSkqh9GeNlS/p7qtmLSv/FOwQbCekxIciAI2d0ASduE8beGuHfAKMzIEPGN9/FOLLCe2Zw
cz5M0seOnokpsGQDzBHJkskKLiQUBgV9YvS9ONGVqXif2XNtvbt7MTDudgvbY2DX07a2udmGedEz
OBWFlN9yrJrP3fG6KoQhUzyOwnM3Ln+bmsUVNlbtpzVjwvkrBbdtGLSHHMS1JZg+p2qK59eMg+oK
zKiKVPEIz3UZuR6H98EZHlKDxgcIH1DrCfEU9GSocZL2roQdF5i9TkMWhe22yB7J9bGSBpL7xM5t
w6TO+dAjRHfxZOC16k2US5FXCT/yJ7fbKDLP3PT1+36acz0qk71cgrSglNhoAj7qyVM+mESlaIEi
Nw1r76P3vBu6CLu0UHXlsuwWPbKnAD+Wl8ldK2l9ZkK0FBBdWeU8huYfAFWpAjInHOVZU/UmO8uo
PB4KF/YKwe7jtL4JbNZNUHiH1tbThx53aIVlQ6KUe+A96TMS8voKck4w5BNzg+q7UBMlPPaDFOX2
19b389U5jmKx4hdJbii+2vSvC67WEVUgcym1mxgsZhTz3Q7VW2fD7ZHk2FgbLYdFoPl7TL1aDs/D
HJ1fzEElh6UWzn0QxdqF95WF0/3Pw21yZx1I4hw7J40KcdovYbdvKAMKmZQOCvsDD5ceWApF+Lox
na+DiSZCkfsu6Ut30REqKz+r/SxpvO0rQG71OdtN28OYHTe0+1YMCBPNwujopbzLPunU+Wwrr2wS
gsfgnal6C2QACnodXNQOwQT3mfB+jJjw7DZ5ogCmNdiDCUYYMNv66Vn7W0puxx6QAGfMNE9Qm5wQ
/N907vAwSCU9gVppeFKLX8UBrYbu9EEyTU3Voo4nqtM/LkxyZGDstFPf5LOtT9woGf82oyDzClDv
z2aMdDsdYqwmzLtXVcs2/7Ah8HZP7UP3sO0eJ2PnRI2X594pB1kG3e+5Edg9Lb+/yxV35F7z8a67
Pib1IBlVIuXTJFaCnwaZRqDu3C68pUGW0o7FhOpn55p50ApOoXvl3GPsPWmXXbm2E7YYtQd5rq/X
M+4NWGQq8VTzEUrTZzTrTaq6r2x/0kwCD3LwIN0RMbuay6aMdLf+jbAVU3eqv2uOPPQh1hV6mILt
Dms38q6ycXkGJSUm9PpvWT0qfD0G3ZzOHtemzzW9sUUNTHT3nqhz6G6XoTdtqn6EB42y9VKiLfd+
tzqqNkesztI4GDiRCBNupfJvrlfeZvZ7vDD4PaOpnhGmkKOjsCThKXN7hqsNFEV/fRUGTYEsEJDn
BUOv3NOcIdb8IQTpB/wS83lMntQvlIdL/wNnq5tBtXu5FXgFVVfQ96EMLClAd8iDt0036fM/shoE
CFIWCEHwvWH6l173voMFVp9yRASRtBVXZzPk+CD2Q6WR672+5rRgBuuoqeWhehyXfgBEfilX/9Of
KNEZgUPQiliVeOYvjnqOgDOT5lMPs5NuTtxmzaPJv3JDvzOvhvwlsw60TUGBRoDoFWJl1RWD3Jhe
qP3LSALBYFdjrih38nUho09X2Yxf75AIS4WwkCteW1RFnC8mAdXTquCdj1c4CPiMj07TSDIBVlTj
5lxSicr7s/0o9ryiPilDQ0p+5W98dSs3qVWPx4tQTVHtG+qBh8T3ZXzx9Vvxe+JlpnrUqTlGKXUS
u55uUS68Z5JE++2WJjoAuMZSyTkxpkBIh7owtGFzIMLMrmVLua8XMMPQkF2AuqiMxz03xmR9LRfM
33482N3dXlJmKyKWQjxAkSHnB7KTeg9MU8bFv3jtQ0IrVcMQY2bxHfaiqaLgmar/uobUL0yFaV/b
JRtcqm/Mg8U2c5BWfmW9bA0l9Xsr8yGGV/cKJAGI1logZTZrG5IvVd1o6os4vIPfZJ5411GZbu6h
Pa5fq+G/INg1IjpH1a1VoN/nECfLdSMinIe+ikhyqQg0q6LdQ9o9tLipTnqgxLGRN9T7RdJ3G0OG
Gk/iuPFmiUt203e730iUZUQxq8Vc+Bm22fPBhJQw99H+7wAmPCthHPhwPfZokfqfC2LYBtRdnxbT
yipujYFB84we6yy7H7Pkop9uFO0p+iW4en197iZMdjYz9huI29dYZuOLdMFg4u2XV7YFkAtCOtkg
U3KyWDGspGnMQhDKZXkbXThB/ZaGM6+YQWBgTXFbFHnE7bEs9Z0Lj1NkJ53o9EQxJYmJp3jpm8X2
KZtVx4EVgEW5v/9fRR9r8e0v9GgS7TsmqAwnr2tK4Jd/j4FE0N7NU0qjmRGxxEO2EXjPf/OEga1k
ZtlqfdprKBobT4rEbcEOMs4mEZgY10K4JnhGsS+AlIGqP2j/i/9pmYKo4BJgZYKLltPHK1n55XfW
yiyl1h8EVMVJcfNGhQUWWOtEq1Ma98OnsA266x3SPcmInjx4lmrcnubqCv9qMJ66/JY2soACzZL4
F2Yz39R4Lr5fLd62KAKWcSOlzi8fHUYzeUVt22hWE1tRxkCCATQXEVAUxjpgPIecuuFPGQICpPX4
Er5qKSKs0jzQamohj9ogHQrl8Bq0fhJLOFO2pYi4iNnFkL7HC+4XGLtb1G6C67/CtJ7MGy216NoK
yfPCM+YaMJxloR28wc3C4wELXF4F1EQdRjasN8fYx5W7xzG845azpbYc6FvYklB9K0CJDWVqVzpj
B595EbaoqH30rFmLiAcJJA9b1nHVNEtxRMIFkFIWd7jiqGw5ciyvkzDZZ4dyGTxOOrm1lk4JRITp
Q5mjcTrqYNJ7bdTsPaNx0WV55+dq3kMyYVUpE5QjT0ET9n9SJepsGyR9qBzUT1ircM6ycgs26Z6i
2sLu56MeSl5MY7nv+nu4jMTPSodp0hJLC5Qc2K/ITnlzyUCh30RTL2CZIlcWNUHOSs4IMNKO37xn
wNlHEfDmpiNqtfORopDuGhBcCui5hb4htkauJYjd/6qMTdLbRymEYtRWk9qqNZMJSeLX+2s+PPoR
R1ysgVLGWzduw/Q0y+V+7kJd1HpcNLRqfxe9oW7CDuM0vDl7OrrFZ6TYW32/PHElQZEkScogCTXv
nvdIr4KMZ1osUA7/Sdcze2aXH/fDt9AuBdn/aAHK7iY9Zr4Em06xZ7d0rnv6eyUQxHnRrvvMWk5G
+JnJ33XjCa60MuT+GmPIrPs8gNdL0CKDjt1s8Zs4weJQgSTa4ABhw30e+YQuz3uL0EJfEcT69+IC
Xgqjv31+7ZYJ6pBBmBY1IDSlqqX/UeJ3JcBIIeWVR58gw5g5mTmojcpX4pIH9P8X/UVjTcGOK8f+
5CaR3x+mH4d3qv0GqOJyRu8Nhd1wJSTTMBQgNcYAM04WI/TN4RuL/cOsYmmuSEfws/phmLg4l5TN
rZC+/xANtZpL/f1N2M8C/OOvIy4JhPNYn2SB1qjMC5bBqlIZFQXcnx7qQ8duVzJli2ZBdFoQnneS
61nxm5RA1xPBl4c1GonXGHlCE3hfQNiigHdmklSU+Bf8JSUnZLEZlviDu/t0GnSO+aev0GlY3bZ9
tuU8igM9F1ZAk7waFr+H+fZGHcbqb5zhzSuDmej+lk7216MEdzphx0DL0JnIoBneTMtdcH2d843v
8b07k1Z8XOmDGEVG+qbH8iwlZaHkJLxokwIiKNLf18ZKqZqCkVTB+3ccYjo9KXQc/Wwu58s3Cq4P
KF4MOXFPQifIad9PZVavsnsR+qhBL+wmK0Zwwc5TzJhbLlUyICPUEvbRETNhFI9CiqhA1yeTNrIP
vDriI1dOaig+BSCKauvNzqol1CUEjwXurpqmmmTipCBGkakIwMKf59DAUa+Zo6KFwYJPpjNLgb+I
/r5yryTky0h2kWXzqAXc/hLF8eTHLRfD8nlvCIL+u5RUXTSfzEqlvG67+IQYrakXOqWL5p09vWPA
NP7bJo/9yw543FZ53/yd3HQRYe5kyVpmhnjajK2sPLiwRMRHcZ7eRjkdvC9frMcRO1V/bo3hfJjL
pnNnvSV7sj4wJaCI3fLXXsKua4lVKeDsxd5ieKwvKE6E6oViZ90iH1d/Cm44kIy8kilr9hqIWmMF
uOBYxRe/SmvjyyWuo7N0k1R/9um60+znT+3koD8rFp7PZq6ZAV7Jav0CLmokk6S6YyX8i/jAWUoC
kVyOvQdtOupZ06KwytB0GTN0jrKgxnBJC10WBZdLqp4vilypFYAgp70CNYj4OItGWzWJ7uWaYIYk
W+ni0WYHOnv80BGAognyStW2aIVy1DQW9Jr4waoKzhN9xuBjnFeXF0jq034WpGyh2kSnlFXCm+3a
xloH3HrLQ+vwrLcWX6MboE5+F488YiPMLR3lVqTssqXeTH8xAtw6Jaw7isajHTljLOoPFRYNuVqS
5Gb0ITOPc2gVe+QqrE2dtddsTsBq8opw5BCbJ9SxiJ+of9f934u8DQFvuedlrzyJxebDIF1nou4m
BC72t2PV8RR3/15Ty4VaZR8KrC/o9oP2vWfy8MnFyYLxYS7/qgypU7EBeuAB+ZQewpPFjzKRAEUj
aLON5+gIlGlrQ98/FE7P5wqTqrqsKo7RPTry5bEjirmXMjRRJ1RaLKObDuRY5VR1j3ADFgc6mPJI
ljjVw7lTQ9BKOClm/D3l79Fb9EztDiSOH8pK4yEc0WaV1JrLN/0Iv58crgNsqjIrHt1autYCdsUE
PJxmd6X9g53Oa1ht0lUIOJn81DU+7UBsy9UgFwwSJwZnOdFOzwJFCVnwYpDVqjIvUR8RATXY9+Ur
tYhdyzxTbh2j0aAh4/rZLsoMQgMKyi4aJYN8U/Pc7Q/dW0/GhOkt27WQMe5ivkPOgHyuerF/FkGM
nExEA0NiN4T0b+x5Vrg1ggpLpDhnvWfrednnPfFg6P1PLkLmmiIMF2dF3cKJFcVl9CFLkspVm1Fn
EDH03QyYjFL4zoXpLe2loQ4HGBZs0Bxkzh4a+imlPJNxQnwfShT6OHs5sXKX6nfnYU4RmMDdhEuP
X6/FpAvjwyEpDFrSZ1rghgHialYMH2SnLRV1j7or26zvXjo+HzVuKuermK/pIdzF4dRCea1Q07H2
iGgDm8DmzqdvMzOBijSF0g+27JaZo/lQkqTwx13a/u69uoPoZmpX6ekNUn2vK5VEh6Qusu0Nj/by
IPdjZyBBs7uqx6+oSbpQDKsV22af85K2eznCqpC1Gs2zim9QLs9mXhtyIEkgnfs/QYgOebP5RnrY
uP806zK+ebD6udUYkg0nN/xXXo0jWRtiHLxKFbqjooxZMsh0EjBy1C6qZueRlu1krnqszgtkknv8
qoNv7rMXHWJaDto144CM0f56tDpdAHfQAmhPsbVxbjAhk/nn3VPpkaNKE1ZP5gYGABbOlH2zCFaX
2a1i/hzwh9iLIHMenWk/RXoIfl94qDgE8k5kUCnrwc0PmXqmhmH4Wp9IMSdVw5O0H0hE1gworYls
2pcSpnOKS2FC5YbKRwtbt9zJrO8oCraV0ud8Rt+1py5auBzNYjxL9xMDIJPe2IXcLMBI1YJrAgqO
t4a3eCU20hUjlONoH6HD+/lcyP+zGwzpQS+Yj8VfzMSulWW3/Q5Ea6Y65Z04I0rmdXMneEAHVbRR
XdQDHN4ySeeIAJpZXi0Y+71iv8yBlBRuNXaF/ispiVmQv7I0sPyLmIip7KxIydJbGvKbHt7tIJRA
xSwI/aAtfYv63Ka7riUnM812El/aosDN4G8qaA01LPrDaqRtS2smpCKaIuKAH+EaEoWhydfBda0P
Fx9XP2Ih8E2RsE6axdPcjSvcjCIRF/wO7bo8+t+vD97eECBo0Bseict7kqx3owxaMhroRwTN0WcQ
/FugCEq6rsWSp0sANCTspXud2Nm0Fxp3wpre0tgVmKE1nvoHliGMR9eaUM6kdg8Hy/QeVGcft7SE
KrBAZxZUSp/PPlHgFvjcAVEybJz67Sjrglqz/eKvRjAcDqxHPI9qWsrN8fJzNsHd+ux458STo62d
H5D+DgeGyqgkaR3CjJyJMLAMoY/P3J4hWLYIVdqkqGa3WmUEnYAL7QZKvHuc9LvctbKkqHJpyknH
Tzo8vsVe6aNffdFK9jwDjcy1PpGb2m6JNuoal146zKQF6nWZUanodbcxJUyggjrTNv0XePkseeVQ
hxgs6XMqM3lnASp2FdTM+l9p8VkyoDBjcIXd5jVWarvcrPan1Hvjva4n2aHlWPwtaIxAgxkZD3X7
Dv5bP8UUqqP97AEo7bmA5vqAgR7Eb6W8Qlu0uif4souIFiiETBzeVVxoSn8EhDYuQq9UCUoWZgLw
9Jp3Z6FLIRWO8AO/eNLPRV+ftAiLlZ/IlltmJeIKgh6BKippODzEIqaBY/bxoWU2pOSY4H81KHSF
5Kk2R/e7MjolQdgidnt+EB7RZzg68+VqqtOVp6TdlHi674DhIbto9cBkeVnBvhbF3thjjHamV/Xg
sNH/holJ56rVQfYxweclzAswutenWCyWt/46gKgEaR/PPoY/GK5M+7kIkRqXf9EOXsM8Z3tQG+V2
Mpc+r8DE6o1MuzZ46fqxT6dw00BdSNzjkPijUipPj/8YCpMkFhbn7RKLLs1mfdIjDoMKF7r99g0e
5JV6S9CcMLosGVBvsueydaz3BBMLr6ApkVa9XY1TkvmdcLmGClTz1IWpDpY0mxSrrJgotTVG97C6
iXzCc8/mZmRMEgjn0Oxp2L+iotT7HD7SDHu6D3sJPdhbWxVH2DTt1O93MN5FCZEgO33l+qLoYcb8
14bmkZf21Hz8tPQkcRiX6+7VMi3/lCJ3MwFoi+pzTH1hDcahn6HRgvmA4uYOnqjGJNnMqomuLw6j
DlQ3wr+9Wd4Px/sS+/+sJ/ZbKDQYJqgLvEc3j2+oF+5TxoEEzB7NIdJm0ZVanp/o9Zi8R2woQiV9
TIumvqOUEs1928w4yB+Tuasu60FF4wv/TzRaQEnhPTcURdfXS0OhNQrEENnyvK5twMoFzyTgdMCt
t4kTemnfmkhfDffKzO8bp67MWeFlgWkqdUslUlXLYJs1GgYwHEF3nljle0xjC/IGVbkXXpUPmEdY
IRef7Tzb/YBxzEbsf5m1OrCI/pmLN3/RyWt4dZWBtsUYAnuDzOocFkx6FCLcVwWzqywYVH3CMtHD
AaZjohuuilAvudC5SeQjPcLs0M2+FjyriKkqYomAyoqe6q37fGM5Z5rEgrRWM20NRIblYSqvBvTy
DKsl4eOijoWwrAIBYbwzhj3zo7HWOjj/iQ8cbCQZuXzOcdPde5YelbJxOMbj++/inP7RU4Jap1hN
kLsN8O0kYk26tdOecT+rZ9ib3tZjdidP7YDmobYL2GA8nCjwLEpANg7aZRFgje+YYQZ6f9d5Ovvq
xUjSaRTsbz7svUzNjkxtKlevNndaqadHloMOsiAW6yyCN5Q7LEAojXWXXVIGcdXTQ4qJIj0a7QVx
dGOuePMDu3MDf/Q2fah6tkx6dseKfUAwEhuau4oQoMuavTt1IoNMMb+Q2BFyi+P3C0fWVwtVqvxr
ipK/f06uyNnfNtfzWdyDAVmOhchfFmfqYd1lq0q1zP914YCKEGP/+/wh1o3mcRsXJf9SSDK/auJm
w/wI5fH/7Zl6TgzKjLIFy5n1SXuhxKCfnbu72GAM8WqfqvZFYlsRhVNVm3fGKi7tG+eyMO0lB1dl
b5NJwiuaLZyiDpLM7Ht8bu+09KeiZ3iYtyVY6V/CdfI4aZO6rSBu7lxejvJTSs1jFKFkuvx5XXRS
doR12Qm8gvLS5taOkyDyAKzJh5PG1RydIYHCHp6J5sOMqbt40OqDKNiYcyxWd2hUQ45ViFnoX+CO
eM+Pd6Kn+fpoCq/IlnmFtYVxIABQef0t8ONOqFZQqwY89DnraOWqJ00wWhCv3FV9EvDiDiRFgRbq
03QFi1HNj+eP52QHNDLnF7MpyjeIGzo9Db2vJF345I2PjscIuJpTIJqAiSgkgoMVqTyVjWcHNsAz
3Gq/ZIqfg9NkNa4bpq40Tgs/bGiBlHFVN2q53iiwoghQJH50D3d56eSw2lnU20U3FAjY9cHZI9xv
u2VCS9rUG+o01CKxvHdQ5rGT2k9aSYn/DlILgwZdZGOMl8BUVKQjENF01e+zfD2Xqh4Eq2hbls8y
jytx6wtvxGTO8gwEd1iKHdmKRmLMJgwqNg3HXKy4SPLlyc00eOFUXndKAnuC/ndVBdjkNLTfnq1T
tN2oCwV+Gpr3lPI8C9+xhe2B8F2HyihT18TGezebGQgmF2rczohE2qlgJpf8VpkUuO4MeKoDgEcY
arx8eyMGR4JWLcPnO/qwsq8LF8KtrXZaXwqm3KRJWI7qGTGK8uYbbzbBpEfdIHeirqU39RWjQEQH
q0s3cSq3a2ZSZJgLSY8WCNY3CenUgqdsIwQBpY+QnFpsYhyIO5rsWiVo5VKogw3V1ZXgZ6sKY9rZ
PpH5V+uR9mgAUWJndQ93RUV9lbmq5Gd8fcpnKWMN2nZ82Q92lzExmJyCMiJA0b/4bWytnhxiWveW
fLc1jYiTl9KUgtvOJZ8utAjlaZXqrCINsXjnQ/+eKNTR7NNtqXZVxWNRInnO2E0/+w5V97dMI9AL
jAD15kir7qSUXqHlNbRxI8+vFyPp+NrL1wAsB1SGGQ9igFSDy+BfRwjqiBJYAC8JKKUTvlsivwPf
Wr1VuTjkBJ0mHUanITn+v3fXq8WbdQ2UR/TZmWkuvo3EMwWoxnPX3VY++7TqWek80DMWC9ZtwoB7
bdvXXqjfPysRok5cO1Xe6uaK9utcj1mmGUzNssihbfigv3xuDEtVIcnxDFoMTds0hJk7wgT7251T
ci1TDedHnIQ5O77E0F46iv2i1tjS7pZBrCnMmDn1Eg2KbbDEIzCFULu/ZGOQfNT5bups0DHZKmwV
8POreITT0ukS85Mu5IW24++Bt9z/b7sLkMv6PRuo3mfVeNNplUk9VQurMPAx+kRVpskmgqHSMX12
zCtsCQJy0McHUIuxJuIfV5H98ug7FsJDXGBjOPaM+zTDKDixzUVPh840PfTgqynjpvNXf3Dg9QIv
gNwEu5F2HWeftO7BNzQTTRLTH4/Rw/RzGQvsuYoMGAwPXBmuHhlH1S4IIW7d+LIzzNQV/5qAnH/3
A7yqMFLq6dz2K5tKflqkxAQJfXppI9xFmnwq8SbP8wy9HNmSIST12t4CUjyb3ISzhZpR8vFDsLFj
CPAzshP5J6e7SDR42lpy4/NdEaV2C8u139hC0TADX/p3I2mYrkpJ+qhZTrpidHo0kpu0oQ5s7bFC
o3IYdp5MUqX0KuP3/GodY1yIivK7Ay+QOF3Ifs8xwBTCSB0N0q3RgNJZ1IkghPnVM2pV6mxIhK9V
LSLTif97YR5ADP9EKtFPwbBAEpL3dHnQ8GaFMDMHIFpSFu4E9xzxN+33SpLyIbHyFIltbU5ktBO1
woDwpEgarA1w6aPX61JvYowhdnPPfgAxEgt3f66q7KsHYSYJ9NG/g8mgNcoK6FWj37UKgsYTgaaQ
r/3mUJtQloxVaOpdv3qFmkEpT/zsHWd2xozHfqRAT8Z9r14ydXG7DEbpfdAlYuXl8ZHfquzedCbz
SuWtKLyefdLof1F0dqoKCfDFoFeTfk69jd39xCnpN5J7HL7Hjiw2b1GaKzIu94nKBzNzJW1+rbR+
wQFvlZrn1tCxXEJlWdl5OekAhiPxPhtfrNzFyWql8nrd9bXE4XPGgaBbIjeru3O+ZLkd16EMAkQv
xT7OQJdhyjajBxe0bkKJZW0YkqyMLU59PZYM1layea1vQ2xmHcXds0LdzY5KRluzaZmz+6lXLygW
ZPMPydlIzP7/S2kzsNHJM1+0a+b2Nuin2EdaaL0YcGzAo6TbQ/M0ajlBGx0f3da2z/vDWZUwZoFm
SxHKPpGAZ5/ZqkM19whkedmPmraskGauT222jE0/mgXgnUHANAcmX//sfHONYMlh4yWMGrDx2DUh
30HsF1DgbaUPUoI7y2Rat67CBM5mpqE8/MZK6IopMWhwkB+NiJPMkFams+HRMEiOx4xBFX3F0Z+w
tVtvv4Cx+nWFzez1TXz7haV/fupRbfNVc2LLP58IXnO3SdFK3PNstGheUuxQh4whkVZINSL4+uyQ
ZEWTgF53Ehfz2Fvn067ROG4GTxF+huUXNJiuWOIMZnWNbxtF2tG/duges60hKija1L60Ubng0wI7
ywWaNxVKn5+gsi8S1hFoVlnOy1QJiXtYKcLTGD4HTyRxBgrkk0m8E5mHuoDafeCNnZ/KV094aPEA
JgCIOLpJ086MnqI4lAI38POgIoupiYlLg/H2GD2OIrGtvf8r9xykPfamxlqHBwtSS3PNnwqugJeI
8ku+5F2UrkYxldEh0+HYTImCk4gEhHqPrPvYnbzlpRHSqD5IdT2XTOHHQeE72mcFYhlRgpj+9h3N
54OOk+9tNYHPU9w4o/qFfycz/Iv2CPPNK4hE8L4xcnbQdbWuJVCM810eW7F4M0ux0b+GUbm8FP8f
TFm7eHLUTMngXPn9TkGGs8zdZIb2951TLHizZf+HJyY1jYKES4v1ogihH2Zo5+r14o29hPzvhXLr
jkp5ur1j1K1JL7eyOJIM/IJuLrrfxBSwfFGt0Uz/vhJOF1vz8OXSiALVBTA/EgC5B4ZTMPCtU5Ag
3jRSGcfhWv+mkpZqvYKKPn1tw+Lp8bNFrs3ZMR1BYtMSTYSIbv3m3Q5+vuzc+SvhF09LAbQrgRTB
L/PxtRRVi9WYZnKQrjQlOIukmVsL/FYjaapv6RxJT+feKdYhjF7E4KymFqSRdaSv06UgxGnq4bFW
Z1lrVl3SPUt0JvbjYAod60QKYAym+XEoq8QwX5WzLP7sVWhKe4MILO6fvSER7mypQ6SnlLfdjNHr
CG2D49efOW9XkQfEU55g2D1fYfn/LVnLR1g3AEI6MPiYc85Iq+qcqXBJpTkWq/bDUT/kUoxy+que
y794DP7HykN8GFcO7YVVkGufQzGCd3MeX6ulMNdM8ThXdOhBIRvHnyIYzTZSOfcoamkIONj9O2aJ
AFKYw58HQUxblpkly/tg0Ez2MLj/GleFat6ka2RRC90PX0CY7Q2AOiUJ6+DbCKYiCKceZqTm+EdC
SF+tMPGC6uwgUb9vh9/VsCeswYGdRYjhyt6NJmK+mwBYdJj9MNWp3YAVUPh7tw6SLi/5ej3NUu/D
Z5P46u1oe2txjRP3jvUTB6EwNWhHnKNGUXBdW380QxPjlqYr/UCLFHoANsujzbIIkazoq9NTuveH
Q18Ai8GQGpAtJ+fvqCpiHO6oA2ghtvIQBBA6A7A5oZ8Cpv9rpib2hdIU3FnUR00Q8Z7HniC0DxEK
hOaEiNCqOHQXHodZm0jaquHothWhodQPKdPmq0PBPt0x1yARLdE5GQyJ+o0T2SP/aj6Yb8zcaso+
qoDEnZt8ncDu2GCGvxf1ekwjlpjcs+3bAE4PR7ftGIeioSCAoaj38gFSbxvG8gsajXNtFX0e6lsc
8PGIztGqHriDWjI4Ep09T0nOlb1gIHoqhv0Q3mYCWqXSBFVfnkCxY0Z0kUmclH0cL/jkp8+PU/yJ
3FZyn3ULy6SJJ9Lqow/xOfnZDshmwozVEh2oLyojQV0ViyLXpSGoUzbhIfczSjOX59rzYop7fHnh
3zK1vv6HP8pD/4ZC45HA/y9HqLoNQDl1oj+UJ7K9btcRiN/Cwf0vjHrq9e/KATjnyC3B8QuFlupZ
yhiE/aKT5FxSNvJgfO1vlflL9zQ9/OVjMe84xtlJfFN7n4RqP523FpYYc7+q7O+VgBpDIEBEqjdZ
70B5edPpZXHqjrGtJVMNiVkccuOYGZcbDmAwPF2cx7keXOR5sJnTI2+CXpPndDuaZ6UJC3qDTUL9
X4FgifzgmKJuE2Ui8NTwZus3SwtQaaWcyfX4S95FU/dpRV4GuDazsaREGBzjqv10lBgkQpNIR8ug
/P90KsvawNX9NdUVyTbwtnliG5g/rXUFyTMOnuZYOk9BxkmOvQjwjkIjDhVSxlnNY0WfqXmSpCFG
SgS1xggYxdVG/jyqTVeqn6Y0z8d2TplhThYt8AZNWknikHie0n0B2rihH/fRRhhwc5jlwHvx2saq
t/WNmrvncatFzL0MPxnfCEISx2xA4CbcTKyMm3dv6dcmhvU+8S7j0tyx4SGCIOrhzd1DToyYbeqQ
JjSoG4Yu7b+ycaUT4nt1eGuJUZjwwB1hm1iayxZyx8Fn/1VokOz1L1THBpJ6fPSAdhpUqPhOtkpA
aF5FNXuSeEJfhupib2e/u5LzC4X2xADeaMAHy5NhpIvUkDZf3QlDQSesS5W5hOBOVIH+wnQSZ4oy
GHKtCRl1PO4LD3kexhhdJIY4ixCc3Hk68tWl0fSyVo342bmaEaDc4QtvK8MceM0UovcwTOcgW9Gv
6v4uryPo+aZb/OsZ6iFDDTzeIMkzqdvswFRkXjBcZWj/S6ppOBC+eisD7CyrAhgOpgVNIqSLXVwb
pTnPavPChFC93b1c3sNLrCleEilcryklutE18r/R/3Ykj+vGrQaeBFn6BJAYE1ssT44cnTa2/sax
4R9oDftSXffbsOYsSPCJiYhykZNNdhdCyGXHwjo2CIxPpjD+xt8FrUYuCaJjfq8d0C6AeCMDVw2A
6OquImTH69vBuaHqr12dAd2hSPHYrvlUCoUEv9XOpONLZEq8DX++IR3HdYoxBk9BJn4hQsFi9r+S
RbZrU6AvQyhm2ZhZPy1j6W3w4OcXCjPlU9MSDfOeLzP8IyUSyeqMfOiPi4KZHoQII/TdSVbbvwU0
rkAGpEtcWZWYhdyRSGJOJlBe/ugIeQDJqqM2yRNgZ5dBEjiPUAJQ0KooIsitY+CCBlTcxpOfCrtO
q6YJKJ5FBCCVcSxS64srowmQykSPJ7k8a9aDp90YlMXkGTRTt8Xulf+5PRc1KHMPkxHZ3Je8g8J3
jpzxgt2uHdWnbDAgoMe8FARzgerR+78DLbjvdrVGddQgGplXBWhFiVng5pSEmxjUFjNnO/oaOcml
pekb/HJw1cOxq30Wo5v9m53KQJ2hGSoH+MfnqLFMd9YeWaahdjBl0y7+BYQe/m2g5Ia8Nwx2dAho
eBO4AyvapM0pjsrddTMMdUb55wFPgBHIbEwqNY9twqWFj6sT2gqd/5h4eIlxnoo1QTI/x9pN0ZSv
dcuwNit6OZH657NclUUjU0k71nEyacdmnjGSjlHeYIqJKEWP546I/2XdUDhA69yxqlrlVgw1rcGX
QexiFytA06qhSHn+mLne2i9dYp9EPyHeatBGr2Ye2AWMcV35ciqgYMFz1tEn4gh+T7IQraQdFXbO
ALVb1oZwzrOMU7Jgb7iIOkBKyYDvCtmmUS/c+ePehCy9ffk9UTe9pVWG6L7STGP0eVgLK4CqtCnt
Nke+a2as49y9Vw3BQkgnjED2wVKJCUe325i227COkYT8//eKFxKSs12zYtwFB8WaMb3LahtK1UUR
g/92t+QyTCtss3KyCPK899w6xaHFFpmYIbqSZw3VBRimYZs6NEP5b7F5w9y1GtE+EFaVTCbbz5xK
GLX6bpxYjhg++PFjjeJfr0fDwoHyJNyempUfbrZG2KnBj1dYqiksyP3Z2gDs+LU0y/cCzxGuFFCu
4Z8TEbqUFiAidr0p06BLvrBAh4OP5KFjjnzo2TZB0K90RlYZ813oGzLHReREPZN3QcpBk6wAUP8Y
BGWwN31ojwXVjhlPF9vaFlRqurlV9mBgMzn1Db9P55x/qVUi6CKzqABtsi08RQnnSa+u4VpNBEmF
ResT6owB7e7ri4Id+muPtOsZcUVX+yWLB0GIQ7SvMN0vDI2JOfLhWGItQ+I/p8QZF8u8S0dp6Ldq
2e+59yvnpxUppXD5as73rmm5GBc0zzI8WLIzNq6Q1hslkq7eez3jkhQ3vYlV4bqFdogkeeZF3McY
sPMfCB7hqPqbhV2Ue6n6xBFCjGg0+UscVzNQaCwPgDM3iZmFb3+vJmAQmxvGtzvdj5TLUcqbCIgg
uNIa/ioeIL79YH7fSTQ+zLnRvhLpUJyspgqNqROJCWos1mXG7ajBOih5tzxOz7bXwu2iTMOs4ew2
mHzVUYs0s6aEW421Rx/wisSRsLnLXiU4B+LrejTebdMIPJ9qhZ8sJZ1wbOunUP7x0tfGDCiCLs8e
WvMUjEhBdRPkynnWKCsV+7VghObYqEZPpGlboYJU9kWwbI/DlU9xffyjkJX4bUcKr1Sumk8BSQSc
eFqoj4rDd54z23I4L7bVyyC5iryaobE2ltfAy/grEl1q5F4VKdZGlc0NYgpU3C09fGT7by4gOdLm
xqmT/5ArISnCXoSPhcpLKsngEovfX5HoaRKC37okQ14s+Lqp08HAhmA7yHVk5qryG/RgF4qAdcBz
lpApkWQRh/q6GjcGkC5qRMg/eAUiA79jIvHY7/TTV71kG8z/qMnQG+YjUzMaVQpzW/F3W9W6GgLR
pI+5Y6obfAEq+mt9Qdt8TJFjIzlk/kftvmMWPK0gElvDLi9LURKGmfabYcXGQ19sMpHy0qmXomnl
TvC4K85WQgArexdwKtEO1O/y6dV8VKhzRoLS3uuSBwxc/wdBoCdAtPJwmGGHIzmFlmHr+53g/hHC
PfjGZo2PwWpkH2gpPkxQJbaMxsOYMIbTJC00I2YTbuE+cFu0mz25hGmQOfN0guMlbgLIRqPrvtdq
a5YmSxmZWyQs/dbt4grKtotfCPGcnRYJhDzHQqGaoBAyCcoA+0CM+Jz5MjwkswLFjLeZpCG0gIXi
WL19qFa49QX1jmVN/vf1tyVBK9gGOWarMPRUvU98L37Yp59kRxDY88TF2sWx3mdhsJKL+CnlD2zl
veeBMiuMkLk1ocULcGPf+RbJVcrG292u50yNVZjfehRJZCnvsjWDbkD8/kUOJ3N3a08y+Tx0rXzJ
+cysiLVsEQvpot8pimib+bRUMx/QfFoOgXASK+OBELaLwZChOMGB0YByWQ7r+uTN0FA0rnyWNY+T
8wuq3hfCdMcRB8yT7DNh5GdVitNsPu6GY2nKYX+xid1B/ftyTNMr9sOMp9m4EOSGdToGry/0Rhvs
oVU/H3HTDBu3/97ioqwiSD+OO1sI9uvjyqVosjx/E4ESoVB5L/Fpi+PHZOGsupCmUhfqNE50VDsS
qXo02NBz6IWirr1U7MS6qu9EAo2UNqeOCNfk6ZokeBr6Ry4/j8MT/PwflIsBVTvRRgJRf2VTMB88
coNizK0vuWDdxY4sCO7qZgxCAhrsQ/FrhCNP6QGRBfv8cctXxfnAko8PskQUkjcNf2gElBFA6pCA
jEg5ZnQ1hIzunCZ1S4HmjC8HUPuR2GuDRBlqxoPJuSJbYyfkKUOriH/lkOHmBPBwfGdvYoYu05ba
WiVO82zEgPis7cETehzi8DmLalVORENU2czxSDRQUHVqc9FApb/Ff0UKeN0zxzzP7aaDNmTa0VpB
pMVHAw7sxTnhWtowWckoh0ocs4Y3SlkoHKtvfovFy6LXFaxIdNTD8vX7jcLYLU5T3F0obRXWw7IH
F3ytUBVnIzlQXqkgw+VGNQ5fjQvYOjs6n+cpzvr+Igocvi9zvH7W4DMeR+XGko1XAps0RIiipesK
nqqKcYZUTMOaWHqZKJ6CoDnRfugMnD9mYq0UYBTBJDJFsY0XXBracz4isbvPboiMLHu2opxVDqkC
POJ09JqHcmw8hFY2lox27KSnaEGGo5fDahiUnMWiLjSWA6AnY+agBrKofXwhZDrUgJqmlkzK1fff
N7OFlR7vH6sqW3RjZjHGPDolybzTROISQGZv8z8WcKYrPvT5ORjca+q2vZHCA2JHVkt4+e0Idz5g
gvPiisS8uxGG9ACWWzFTvQCLQTbzXppcgNMSfyRlMN15Xo3+iYX9OtyAn58SO6O7hHgN0HPa8bEd
/IeohdZV7pEZ1DOhAN+pwELUZSXfUgyCJpCvumesvsX5arhwrueomss9Vjmv8XeflXKQ1sV9mbR1
4floZZu84ODdbv29NPsxXJoteAfZnfGS2XVBzZlE7I0hALnsV6bvah95gsxCaxMoxLS/zxYRljXU
MNMrE+s09l0f5v6mI0c+LI/s40xjfcRfxr0aPqGnZCk8z7oaXzH4rO5kBqP+SiY3I3vMgeM2aUQE
1EG3nzwjn2PzhCf/FQKAzSlRleSaYw4CRCqIixRIvVhtAm5h/a4hTLMnvDmVxcfKT6Nq6DTDshgJ
YCaEQcf0xryzc+C0e9/Ll0zGQmU7sNAdr1mYNegbDwmv3RcR9jMsBi2pGl5W+/6tcJ6E4VZLR/lu
ZjHU2cE8iWstU76xT35mtjMZB2jpD/JZujLqvshVpDt7TQHSD2noLjI9olFQVWEohH6QcyBFTJ0n
6ZFR+aMXBiW+baqqIbTBVOwG29qQLXhuco/Ms1TAhFv1XfG+QjEv11MF+ExKDe0P/KvwLUEq+srF
NJ/gWuvgfeB/tU+hfmws9t+b3uTnsVgzgtdNjxCJ5zPpd0K+0Ol/1udddS8khXKKj1EcUcN5dbBM
WNGbQrrp7b82a3ibhAyiZBBNIJ+L4sqaPurnkNm8W4KQmDoTn8aSXFf/lmMGq4XaHiRtkCSB0ouH
c6ZwueJxKHw8x4RL3uYZrR1e1WZ86XrlvJaMxwpPmrCRCEbXrVnumLxRCaE+oNpcWwwy+6E4flVx
gNp2Ds9K1b8rcVNQKFdp81XAKPQY0e8kB5Tjyc7UHuEwNIzZLX+6h+TIdAJ2/xT4VXqhVFc7RAVJ
bQ50fEU3cw1zpe40GZRV3+9qZOczy/ZHiLXbPADKTA2RG6QWpffGjvRmSrzXrho6gAUrXLUWNK6b
4j6S4eBB6HaPk4X7rjS7sVFKZAFGLamA+h/INiD+OcyYc3qS+RVx0da42GIEvFMuj4xCPd/kDnyw
MVlO8SczOISJSLoG7ufmGR5cor1bnBfj2gMdusrujWHpnK/kmARl23sIvBlsXxq/PKiSVAvjf4Yn
MLjQuMl+iAYBJqe99YbFybOWn04cLKYkiJ9SolF/7oBEY/rIHsf1LaVWdtE+QgDN7iuPbRhKndQm
rXLNBYkVYv6qtNg1WCSyUNY99mOo4eFOCBlORP6BOLOtwTjSJONI5jvqtp6DXCssN2nWYS2qte2D
rsJUVJbLqNwO0ZqYU3xYrV1s9WVvN6WTGJZm9rCjWSo39lJodQmSp5ZHtjcmvrVTNDWnhCnTWKzy
acZAoEFg1G+Ct1m9v6rCBxFDjgS+69NwYnzSghJ9RZBcmsIlo7hCtUzGQaGrDlKo5+Umedoq6MLg
J8pDpXukVW/2RuYx6FidSsK07XoLxGhiOR2pWXFl13wB/OaQTVlo+52pCj0mdFj4GwpArR5mLW9t
LNG9B7wOjVnACWXzDW+qYpBxGEoo9yunoS54DOYUd0ZEunSdNpbPsx3SBg96riU6Gib4ny9ZJu8R
yPrXvskPPY8YXWm6idV9k7nRxgjT5LSC68DvMDbexN9tFe/N/LE3s4X2yklGG5vrvRHrZT/Hmv+H
jP1In4q81ZxUdpv/iH+p+dtQY2Pe+8hlRj3TXMLBoltkUNN21tiPigOUJffsTTIYEOfj4KUlMPky
qqF9H5NTdbjOD2uYhtgUhPFVj/Ssq8XBbgbIL2q1Jom/1WTIO4PozjoEi+ka1f9pd/4nA4ssIZD3
PLjMi6Id9nF9QEddgSsAQr0E3v6zWdQl60EV1hK3VQw1VJrgAan6nV2blDRcbTR15UENbssfS4u8
j5NlpukYZBeM6nEXuYkGuJWrqSlriQJPX7loj+OVvN1d0N91jDNvwc6OInCvv8o/CjQQ4sT+WS55
w+bFnpJ59a1qG0yHDwSbhNqbsuMqPqcUbDSYtMtAWfoVwv2/0yidmY6g6sKO8iP/3IndQcqRB6+y
oqZhaYiakRZFLQER062GdtbtZ4lEczLQbvukLOLajf/yDnSOFzZtfUkrA9C+Hyg4O4+bjT2dx49Q
cG/ncibsyXvmwyr4NDFdawdWjqlf3mdOE1rcOTeSGKmqgsTeEMWOVJoGLLMG32Thooa0vhCty+5o
+BxrFQop4Z5/hQ//i38PV+QyiqjP4BBdPTcICquxN9ZqDxP+zjNatspk0N4L5Uocn7SVjYaTZuCL
WQZyJz69fnOYgSLAdphF0S3DKXbNOJVRtaiYksIN1f4Zi4zW+2Z+tUza2kHLj2jYz4WImIFcCOIP
0UN6B0DKI5We/aIWcJrW0aL8z5QZXdrwfCKnK+ZZ7maFsrwy9NDOBbDzxehxXrdHLZ2IOMc3P7nR
QVR36k++2mvh1iFGlSm0d9zbqufnDZ0oNLNmUTU9TcghuBqRRIAnzFRnAY9OWG8vm0C8y7Cnv6wd
lM98gKuO5kVVK0b+vPQiRy0kk9n2YnL2JQs60pL+flEfoPac421EecM/YltMJZb9lUZhHaRuSxwc
fXGbScS2oz20HuXdLB0RS1mtLv4Mez36w/wqjBbZ7VF3GmpYm6Xsp/sg8ccmEOTfencCrW5vKPQM
RheX/UtR449QohZAoNoz/1Od8z55rjx4i3Bli2fYBHEWajSLcXbqugR8s2/JxddHrNTPpHowNxAR
c2T6DyzKBLMSgS6Qrktc2mAZ6UyjGiFYYJkof3SuBt1cDkbxKTCJlLUwq44OQQz3FrgaICyjFmZH
n5TEP/KqjrvcDKqwcYcQGcK/CK8Cw/XSDx+F3RM9pqnbX4FMXumP1BcIXvh5Kiuaz/doE/iq6vMD
yTix0NxzLiYqvp9WmpxFowPrzpHyG5Ysig+RUWn4tEGaa9U2BdFu0qeX5vFo98L/dV7Fsrjke2DS
Ntvww2yk92vSdDGK3PY0WJRodBmFdvLjnVGVoQnT94ohy3/ctikhPyppC4mIrdFamswvDsGBhHPF
V2DT7FBYJvJ4ZBQ94hNHnUoptrPqeLumP+96dAzn+ZCBLkN0Qn2YwKx9eJAbzmFoGIGcyBRtiwJZ
6aAiKDzm+8S04MRjGp/RbahCkB+z4O4cGcvOAwZPuoxDEs94DPzsttRpdxFdYdJPz7kAWdMky+Qw
WCi+Hmhpb5kiMOhrmWb2c/zZb2UZJTjczIhrwYUWq1tGrCilDdZD9XEOC8/1fRfRF8E4W/ZNZDcw
3zslJpyxZgXWei4pwKb6uEjNmCFyYrjgiTFNNbt5kSk6TPrtu8ljS+PaBEcmsq0m0oNTeYogTyS7
8ORYrfsCMS7a4qe6hD7if4/sDY6V2nkNNymFUqspSl43lnPvN075yxogs73t1LOht10bPlQB9rCd
KtT4V0u80WO3gsz0O/OSgGBwgAcIKXZU3VpzQlCAkXg2qBNdgj+t2sryMQ+ZwJXVvH9ELfNSAbG2
lQtPlMXLwROZvL0BOkZJsvS4tBNP6q+Ymc2uUYtNzFT135v0efWkziqgvkUvlsKGULnj3wdLSZ6h
B0eZuyyObky32tyfjitRUFKdK0gOJQNmeFUMwUgXSHQK/LPaMQ195wpazuYsnQ+2XViG7X5uTA5v
hl+l5OYAm0xUGtD9/LVlzvAz2bQsVLI8IPd6sSC9xuxBo1iBnILwnTzFw82wGcfRqD4YaEyv36dS
0kikoTCW6AJABOURK6CRDKZ0h+I3AHtBYv1AxFgkpLXevEhFSq1lrpn5ihKfop2EyZXPR2YsgAzN
GgPCzSSei0HcEL9VHaxP9ruK5C8IBORFUpuIrspGAtZFqLtqVhXHG52PPBMJWeDsLj9PTHOl7nWR
uuKxAfDQwB7rkWX6XACIpXje6IeuCrXF39dJwbrxc7Rqey/O6UXiF+qOFb+BnArD04LlQn4RLhCw
Z660+70RfQgCJy5GnpGRY5zMHf28oU0CFuaV+BjtlkD/6SEKoLdUMZUiYw8KiTzAQemt6eT7w9X7
MuVidSHy9J3OWrxWuzUqSdh64Zsu7wcRauCo2IG5l5owF3/uqah95xb1Md5EQtsKMJAXze2qYk8l
o6Ww6lQQDW2lWkL1XFBoQ6otKYNUNBxCMIGrGVWFe6X8rWpPWn0cKdh2pVhdjTQtw6hu2Yo6mLk6
st+B58zHogLvjMQvohqtMWata1oQwAHY1bZeHG592rJuTxEfu9OrqkkCYO4q3Qo83rTEto55oZa8
J/bjrZPkrBh/fiWL7MdQiHLz0W2sPduRx7jFf65taxN0mCXdrOMHTHSP8qu6PwadOeCLELYC7JAr
u0X49/7llAxjRwm2xVbuYQPUwIudRUWPCYSLU+MJGRBg6hrtz/vytfWtb+rPs4B79gR8gNW2JR6a
DrZT7Iz2C2AcoLu87JwHbNIJHItEGcwymoqaZvNs+t4jl4Bpst3MEKOg03I9Qa0j5ujUyaWdJiIi
/V5yfGoEojvGRQLjbzoOwt2FL4fQUfVkiQhvVr2DVJ9AwFj6o9EreDRI6AlMyV1aB0hUEbvPWnet
Y4U6PWk7fIHlJc1Gd31Adp+vjqJocU2JPYrvBn5u7LPt1Mrw0HH0uMu3F3+C8makIXVPnLrPgboD
K73DIsh9ArU3PK/fWS829wNZjsxvUB+Ty41v4P3uJq5gztvlOdZpu7Ktke6P068NtfjQX42cKn52
F3s3EJBk5KVB3ke2rF4ufBKzbPR2iVKwpnspCNvNLIz9QQ3N4H6cgK2sUw/kro8iGYd7Ms80kmnH
QuN7GuuCkWLX6w4Xq4alYeqBy/i6nAf02rTyvj0O7Zw1OUkALLAu+avAjgUXi2rVz/2EEmJHgTw5
HUwJu5c/6F1zUTxzzXkx0C0JrvNtSx17kpod8NhcfTKVjUZvO1ylMt1/QLcpj+ZHQxQTLuEATIBa
QBL4m/a7/xeUECCDz5gjFNsDx2njG2UPykjDeEjGzNhxl9osy+Bmo/FHhL3E0GCUp2StzqlX2BXM
3RV+U4mKvLFDrJHQp8/G1rmqcuunaEO4JG9TIqAw47YaIrEipTp6xrRsO5+ipdU8l+PQL5A3NZsF
PIlTTCzO5hRXk/NMJazyXoS5VYbvSXveAapRLCvBH3OCAz4f16jAnsSC8zs5eVYcG9Z8byAR0fbw
mDVBAqaZISsUXpYXGPem0+976LtwrfdRGjqY1R7vFHb8itR5kn1fzGXy3AaQKniON0v1AmszuV1t
dzfdLd2/SCb8wzu2HevgoL+poLVR6zzpXKgxiWhUQMZGExEwDHdgwSHsBee7hQR3S4+0zyBAxmGm
X2V1wOaAOQ9PaQ2MV+gSEmMPZ032wQHdQbdk0Zw7zauJHQ0ajgLXSqVhFHl9ZgNdNiq11+VfHW0o
J7f/Cv3HZDnmJX7BMDKTRUwPJEAhJb5LSPC6vmoFvVvyC6QLLXh6/8JSZ8qFQcEsxfH12UgV0tqa
Aa5niLadq371+k0SdqAMpVWpsq/jrZIGU17SO2OziEq6nm8NWMVL1wnzXg6TmU+SC3ODdYw0Dhms
Dat/hnq4B9hDFzURxVhPaB7DirxcvBGZfIYWs5lCJY54HIet0tewxhCGrVBYe0i0lgIZteqedV4X
lsperIa0Jg0EKRqX6qesr5SL4AxXLdJDXhQKJ0HWFvZn36tIXXJhip7SNPCMCMGEBpt7hFa4hPna
DZk6MYYKZ0/uxkjvDynklJjIfvvMs0DJzTL8K7M6nYfYtJR2AutGko+oO8UFiT0f15C8ASNIkb0T
ISH0K1iPk+PUINOhF5QXbHCKMOKCwBFS2IvcYEPRvCEwwZonIL1UOBfg6NiwAyjJqAAZo8q8naRM
BX+uEJGQvIWPuOfzvHHKxexnf+w80HLg4DO424hMHf2GePTWWl646wgfyI1xXq3LZ7Izqd5SbSQT
D+ae78P85LFZEkY45Db7wj7sQjsDeW6TRY8kyQPwb/Yvipi3WxoSiSKuQS3aZW0sltWCtXpm8Ogi
norkzBgkY7zClMYWiu64/tTrIh8s1p4117pum4JTPxy0iCkbz6tx1UAB86VW0yVxLAvo3adUQa0T
ELLNtEfLujLFgMfwD4BkGczJB5BxKlckaI7OQgmGjdy/bJIB9mKUJnf5CEz50AIgAOwuXVuK2G6q
+Qs3ior5cSmdAV3XAs88oK+tWqIN+H2SRBEenI77itV/Bvm2lHfnrMnOF+onEGr8rYxtXS76i1wg
8rOCuL2NbcumzldDCK8uUHYKw11gT7KBK6hTf3WZe71rjrtVacqThewmeP7R8Fov9R6frb/HpZ1z
K0aKV9TnMbDIaBCucLRUVxTg2h4B9wzN37/fCNLpI0ilVJZF7F2YRjVovVfC4xkEhqIQr8uQufXA
ivLxFDF6tvhayF/JUnXvlN5TceLqVcnHeGHq6zeQJiOkgeQe6hToMwjjwz6Pv6StrN2PLepEZM8w
8z1bJIxK9a535oWG1sIepCNpRrMM7i/jn0gbfZ5TslSpPq7pNrGjf3swO+EzytWjYmxwlD0z5f4x
Q0rU5WM/OtBts1jtZMEjglv8PNuDjAVncB12lGzHwvxxWoEMkw6N1j1nxekQ7FuAb9Fgz69XsJ0X
zBHHKy7AB7MdgGonRiBLn9IcZYZh+2KFb7fgS8Qszjl6fdfPor7lDW/NWZONSS5hxFliFaVaEE8D
0Y6JUWbOLCMDaKd9P5w9/whUbk4t+uEUlKwNW6sXqwZqaCWeKU0GUwVqGWvgulMvcE7sYuRUURia
X/91DFt3dld8siDJjb+Oao6fs8LUVP6eS6AXY4hz/MIzKsB9WHABjeZ0/D1VXVVz4xLgy6pz6lYv
/xJ7lHgnNhndSQs3u44xPKGng9tUBNT+drQdco5dHA+mf9fvfmEZXbdyPULfgr6dEOBqEkzuk90r
f9RR4D1sXGAuP3YYjdG5OYe5qD+atBTGNG+ZwsjyQpFYSKwxnbd0TZAOtJXElZyRZqBv46IqDVJm
BelW1T71bctsa2MI1vsNsD+u56JBLCkP94HlCW3lSNTtDPsJeUkGQGdfP3PcvAFn4WMmMp0EKsOA
qgQL3AKL6KgVpvUaH/rXECJl94d5TIIVUCgSSh1bXs6GYnjs/EkYDl2FuQlzphm/Og02r1iAVPxS
GwB5UG72wvD8JjjbRjgPiEbOWPXjIPQDA4WV/nVEJC+hFknHlE8fRozou2GkD/O9kDESMsQ30mLW
DNJ7/zFfpUlBQmKf5DR4mUnzWNDo8iCU2RD+x5WeAzwWMYRBq2QYkqUG6zBhG3CVgc7FepcyV0ga
xYiUsxIQUdlgZlkxLqH7FmWiZu9OkKJOPJAgRGuvPKDGG9NwxiaeVzNdvOuT+3BbFkjOuj9UJso/
FXuG+pW6EuskRzdr+qR1jzzv1WANZCQODQ2r8egOh/JOVR48Ahg3F/KrzfISQEj2cDMKYyQsnTK6
PHFBEBLWa+z3Qj3mGNnH236a0+lz5ISMIrJE33kuq7p6kmLT/lZAKM3n3Ldua87L8BOuf3oW007P
3APXkSORuo9nVUvuMGXT5GT04lc2pd8UHV+shX4rOjzsVopLh/aR7pJ77OVAJ7+GBEOHcVcYzdBH
lA+stOJlrwqGqmqCLSHz1I55v/WmNHsvs04ZOzVy/dYBfBhaBpmd+kFh3XAi/haWVgB1M6sKvmz4
XgBvLbNqdVrfWnUBeVGdFKkurC+ACtuRTNiJ9CmDfsOh1kpr+S3Y50VKGzhUN17ojYP6EeoEDbKC
XlJuVYXcPtWtkkTosNA3DN5THpfoBVRIefpTJcCtHAv4SZADvqFiU6Ux1K2ubBwEMLjqu47UbkMg
z9Zgkk9Pwx/uS0V5s9ts54u93W+neruLIKdM0k14WHxlOfu8auc37qFPguNFMQZKftIgZZh3teeZ
HSw/+VFvSVw9xMVV1DXwgt5qdEA8/tI5NG8UMbq+SPZR5/9LnKirhQFRdGzmuMrVegVAJMPNXoRP
K+W56d/DnqJXpWMVDv7s3BF1fn5cS2AHa+ScKwCkmRwNIvGf24/FajTBJWDfs2ZB5GEB4R4gl/rN
FdW98shdiiRnzPiFf0GRb3csOI4a7q9Tlg+Av5nW8FDOpc6PiUV2ikCSxy0gstNqpKCWQUwcSGyk
Pe53iJfCA9KrWtI5G8GGpMjtOXMlLO1LeIa63MCgBG7bc8FjZ5w0KF3+SIsnp4SaMzjFBMvctZLS
lhTZo+BIVe1I28HZ0fbDlVvpcPAYep3Af/GXmctlpPcYZR+XAWzGOuVpHc1QRARrXEqotx3EMI2w
qGjUrMNHgM9eI3zUWJ2ynr5bC/UTXu59RoBX8R0URswPHksvF3fmSpU1fF3omrRF1ANBkeHQpVa6
MpeqIHHwd8lDSAbXX0XGYzE/rmNRRPz5hNAXasip2NqClNyzi1hMGkqNex4xI6qE7vOuyJsxIu4D
M17vi4Ow/9mVmzEKnoL7ctFVwtya8Z5rV00VfGQ6i5Bx7m1vPvHNFXzUOxJVAHaDPgjbS1v7f1p6
YELQ4AvZjYGm5kYII0a2Ujaa9E+bWdifj7ZCzN3VkHXQU+dg53A1LulhpCbjOvhzfkTvwCYfg5HE
ZS41rZXALFVrrOLyBJk0goS3WvX8eaELbyeAk3v0/s+AjQpChuwDEjj1cMZLTWktp/Ii/UgM5Alj
pBzk2NHJKVt1TF7s3va0H1pOUOB2TP1a2acWWERmb1/P+Bt14I2RM09p22rzZ38B7MJGj440O1MN
cdZ7lWR5oK1KzC/bZFc1SkPWuDUSJ3ECRIyOaqp0vs59hfaA3E2Dq0BUthzjmwPH/I9wELgQmKml
/XD187GTWO1T/k6QKB62Zhiq9qxYvMS9tWYvoU9jHcGnb+XcexmzCkbf9FGnP5XWd50IJB60ziCX
U03oi2tQ7dqmyVDBFDQs+RLxBNgrC+iqLmaAA19ZV9ASr7FJK4U+tDUvH7hZpNKUbj97icwTgQGl
yLWOSJOTeqAxv3auNFGPP569WSrAcpmYw9q8MgcQVF8PUl3J7DOu63vEELZjqvLAvZlm3pHV+dDd
oFMnGVuuYHcwDvsHtag55+C1X+0Eb5lu2FkTPwbFxk8iSr9bcIuVaIuSD2nqXRuR4AqyeUhEEOeP
QEFlslS0YeiWV2a5cgbK2XWgzqyQ8ZEWara8l+7xmI1+PJXKJwhZSewMpFnbkM2bgWcJ+aCx6mxl
yT5m5h/WfMS393YcEh28hAFFPZ4TW4gCtkF5pLQwSPNei1DJ933R70JVkag9gymcXnlnViIhenuy
s2x2GWlfxIwQvM16OdIWOYXYFCzMwtH8cuUDFCT37xonuUS/GS9Mf5q156ANNs3YzuNpPU/p7Nkc
v2NkygvouCUzfZsnVnKrX3JXTAxf8U2QlPSbnGmDCzb5KjFcs78rXUguFqaudrgZylLvvqsKQR1B
Wx2beNRjKVz3EQ9mB8klr8Bk0mtZoMnFiE7R9T/ig9kog7GR/u5slSRx6NLsWwjGgYaSWDtry6mX
OkzVEU2FvFQZfWi5Rs5wyWxNj1azHjWDQqvO8xEkVWDqq4cVv1p9F0fsTYcNx++AoIia0OZWsMOk
1UA4v5+MAKKCFmEWRHYJx1fsq+kjcRWCYh6CposlKZsaDvQgQUIEG4JBQYTM41dKEyFGKdAcudpp
kZeaV5H9lrE3Ak815wtuPEgJg/ON/Us/hHKIvo9wtw8ryazNlSIBng7o5CBc686wF7kcaU2bAKD1
uMiCUSLyim/69MYizxBb2E/btjfp9smhlDcekr4Xx3qY5JbkvYuJePyhXHyI2MGrf7x2p06CYMr4
+Vt6rOHY8nEUmpxCx+HyEwFUW+NhmjOkvhDT2wZgUj9IlbUYZVQ930pASr3Y/1sykBFq4VvTXzwc
mK7eHDajcDCGvFAS9QLfn/8qMqGnYCT9NJFc5UCu9T9ahyBqE96+vuaEly1N5nWYE7d+IP9GkiAa
9mUvnjlAiVF0e8YrtEJ18rY8581NNsCZw4Eh1hkdraS0WgFabDSToqzeFABPMVsPkzer+BWBn2Fo
dESgRMKtpBnOK88W4NoWAqk4Eg65tjHAh0IrmiWxzEfWUrbz3ogR7+rBfsmeC1bnt5YR6n2RLz9V
kpGDwWXSNHwHRGhrz41OCTbU7r20xu0XdAdG6uxoM9NXYnZ0FdKalgGR83Y6i2B/j3nve08KKL3E
K1Hnyl77oSQ6lC3gZLGVSDTujWL07PQY3MH6O06t+ht/ptRr4qsRp+G8LQAqjsxLcfQzBwDhLK9S
xwitjwzAEgYrnxNh7oDmpEoIrGiXLMIN7tCY6IRlORuRaaJFbwsRarlZwsDMlSmjQbbZ+fxpqWVx
0pS5yOU2Bcc89g/bpIgab6kqltivhtQXFH4LRt51JLarhzkHX9k+h4Cfz+HumSZ0Jmet3tzk88dL
cMmlFaoIqB0t32l8ETuaif6aQyZFupLc7Jhf5LRljXwVofSbXsMy1l6rY/yvWNtdKNCgPEuGeoxR
/4y3V4CSOFJGsvxPqBh/hp5Gln2vZqdR58wOk2BzeSIh9DiNCigEki/7/4z9+1nKcK01fGBxff/n
OFRiIRY8oxaCUI0iRwX96gJ8GPqcxQ3AY2RevWBFAYnJRppGnP8XiPnWZ/cKLHayTDNpFJMEKU9D
M9kZUYeJBZbP90XoLwGkileEONX4LPUm0fNCOGKoUUjuee0rF3TiGui/q5keVVB720kROhH8hB2r
yDtlAhRYrcPYgv30SpuFlcJao9AwEDD1OiQrRYqNi+O3rBXPJJcILCS93Qy0QbH2EiXQEh7yZhq4
eczM9fYx4E1yub0BMtDwz6bBM7VSBouCXagMrYvKC4TzgMf1sS9N4Jz27fMlv8OrCEhkSGtKdrV4
6naQ6/C+zWHCGkGaqoRQ15J816ejpi3ZgT+5b+DbtYy4QlDcc9MTtE0by1/5pJNkGVb7pwJz6Ho0
/nrPw2fXPiV4GLM3cFN4POSq9JGWcPdJ5pzMIpHCUEwho3tvip3lwwqVRQ9ewRwdDxYj1BytBhSR
ySc1tvNqv95NAYfthB2g5fPUlXpskoPA6p87BSNRn94/H6VAVfcEG/5/CrA/YkmPpTlrKmXtcqgt
J9DQ6eb7KsX78TPctlWO0wRDFEkjWlw7ryQFXoyrb5Gat1oDzJ5Fl/SaQFMo+Cxw2TvRcwnsrIZw
u5fcDjkY095lVLnQohbzb4dDsX4A+qdjjyP8v65SrsMzSb78/w1PfZrSheAFFSaLM7vUpRy944Xe
LDLGYRktL/Faty8kH54DMSXXeZQxDsY4LrtvPEssRHI/8bXiBnVlmnavhIwaEJhiU/jwHQHRQkvZ
6Xza/qtuz7sH7sge/efXiSa+4OBTXEwLYALYlBU9PxYsY1jvoiHkMzbVGAqBITi9rti95SxD3RIF
em1OhQ5LD4B0ymIub3E+wGt0QqauS1G52vPXRRkfM78/ovNW8NgwBcjOq8oCJ1ndOOeGDfMKZFC2
eDZ1WD1AWTOhIVMCjQkAu031W0L+8qDSF1MiLVQGp14z7Reljgv7VFIKMJIqyiBcMXjWDDemuyUy
yN9gFwm+KEP6r2zz0VaZkgaiaU07CTjIKuNCmDiDkmHJt06cO5DtJOHLmHQyux1P0Th98ZDAPxkY
ztU0yctzAqeCq2jvGWGiM3z1/Xtfs/6CiJgEUwBywncmQyS+JBjcj55KHEyCaLcR1glkKAylTbaV
DHih2Tow+Tt+BVCayDe+WdNSNYb9D7ueTQT/08blqwzVr4/TU4D07iiH3Bj0ApmrUmIfAgVwmpJB
5M5se9PErCdyAXl2N9hlaBMQJBO0iycd5vyqIHXwKhXpCVWEAbfxROT+k9tToL7sczgVM75j7fb+
aVUJKuDHhkpVkxBh8tAaGW3gAtSVrxjTsyff0OFNEvJ2ETKGcYBYNpWY1LMnT3lYuXDgVymaixoy
czlD7K1Q1f8hD2GDHA0bhwoQJKMlqPQm9TLQKd/5j9AWfiyFdFh7pVdBN9V5DMUctsqK3o/bm64C
qm/1ymswHAyIDX4aSisTvNbInoxdJVqiw0NMkuxyxYrHmwHu93aJglxLnmLU4SA4LPgn+CjA0pfd
Tv3KQhCGQydjY1qTRAEk3wB12kH+1vd49wKxjA1S8mIhXYCH0//tVhFg5t1d9hSTFM5TaTzbzSGH
aIQW7W0Xl7W13x2diHYNO54VEU4llc5o8xcPZKBL1uDtCxGjxk/QQGzMjUnOWixQYYnhhNjNdYRF
xEoT/cX14ajkWejZJWt54jOKl6Fi3YFQSDRV8fUnLNMMxyulaet1aGwMKgz9ACB4nrqGHA44rFmX
yzsKsjoEtSqVT08KKygF+5yJdVU7RF8+hWxjI27M9g2EZ5gny4PMu864Wbo8JBhB9Wm1QqVFWAnX
z/44vndWW98ndchI88j2gX84fi0M7k543GlJqDQiffQgWETQpNEYvQZpx6pOR72OjJSYR99JNe0r
ZhPiIxl72322Y6WoKOJgxZIcKX2888y5cav4pmuwlEvkn+Oq1TYm/PrWyeXK3S8RfVEUJDph705L
lvCiLR9XTDT6P5YhrdGcFxqksN/qxz37Y3phcqtQboFpF00uXyRQ3ilooIkNElwN/9H50cVKr3q2
NbT2fc5oK5Cf8vYy/lYhVOXlxUQKDRfHbmFowvH+Sr8PqVXJq/0EB1sGydWQa1ithD06mtOfqiyB
EQVDMyokACbxmUdZRVKcLGkfq8kYV6ONdvQzg5FdxvtxGgEsESISecat2f3h99kDyJS5GqVF6uuV
paBnMeZmp0Qpbo3rgisormWn1tI2zIU3VT2trN1vWK4gzYhPQmN2avjrU1LWBWZ3f1e3eQ2DSJPV
ILDh7V37qgPN9numdOAhxr6URMvOJrmGnLOm3zOjYGBzUlcOtO48JP76QshAs+UYVMp84i6asyai
dUU942LM3CCHyMzhyXI2lnndN5LEtOhw3ZSd4nIhxE3f9Kamxuba/q06FYnhX1GhjGTNEEdhCB+x
TpsrzLwKN9EpMaj3KWdOnh6kbZF4/ouJHERp+y3ORrDgMu9lMUhfelsiMEU2cy77FD6OQX+QKF48
5YtfI6b++sQHS2Otpzi75gSbMMrGZyA3MvDy5GFG9oQFXG7ryN8ZcPy6Xd6gYYRg2yyb3flTVJiE
VR2a4q4Un36Iepdo6zCi07hC88XQBk5hHNnKci2xyxBJboP+H2IG022nTIjzJN1WITfI2zYkaXYX
p1CU/J1qtLbN5GTxYLuj1j1AvbxDAai0r7LR9QnAYikBuYSzGWPm9k+efEw0/tt06MuG+TvHjdx8
BOpkcvqowxOkL9QHVt1gIYouIseUqA1H1rOL52kvXlPnpBml793ehc1Qq1hxv+4GO9tgm9J559f4
SqKq0dfQClZbynYkvdLBb2ouqhCSpCSCYERgJO6Bzl1nPnpLK+bOpudyHm6LrspI/oZC+PbRnIrp
iCbvx5RPI/ITGbZn1lLUcAb9xNZV5NcWYELS5ffC4AcspDECeJvfLOgC6ehQu4edqYWsF0d03SEU
IYzbq1AvRwcXicn3NyOpMlNGO9SWlo714zPfkOFYoZbIsDjVGFwCBeuVoyG81t+17s+3ftaY8Q6C
33Mf7GowTtLs/Qylb063KZeXPI8B1WJds1vWzFw+dKbf4G0ekS296YOE6BWizx6g/YuM4pHDtjQe
cY4eWVDISGBHTdgJ+/RT5Ie5qq4KRGrjSxkQ8Gk/z/FepBmL3G86rzY0/hlknsRDi4v+2tEmcOet
Z2UObX4PeAlXpn9fN00WQjE9yvGQJkeSJHqxJbEICMTDfcogvkTwYf/ya2Lb78WeRFYrRdkofT20
/IjUm7Vcekao3ZHnS5f0//wx4kN5RL3HCr6LaOT3sRlf7ymEAb0PHa2yXwsL41pffcHH5H3jNx9x
cQhYGzBke6RJLZRsYeo/CJcgVJSE7nAxHY323eoRKbMNqHgkm+sxjcHz3qfta0sHAy91ego44H03
xaw3gT8Wj1h54eAyp41jVHYzFoVN1/NRdm6p0kAFiK9x6maQ1MOgxdDkZCHEf0PYSTf70cxZN0BG
qWlhATLqX0GEnbidVyakh8YbLYVFTDKfoUhMHLz3yyJhwvqmRRg1q9OWN80JT9myjLerbUEjq3Q5
uLVylc76iWe6JB7Agf/8AXNGRidNOuPsNRqz/y7Oz2WzvRCtZ3311o8rB388/lHfSeTy/nwocrdN
NoWn1gd5fBR/35mln2277oYjyLCfFxsdp+CwWzIeXTHMj3b4p1IrmWVCCZ75qQYRMWbOaGCMX3nF
/Q9eBnMj373bCHCDuHF+EjbBBBuML9LVbhGhO+8m11Fx//038joIvphSZNgAAK70j2KAXRv7MTew
xtgxseo8mgiQzGLHCR0+xOBIp9Q1KnIOquIwuUXbYUMoB3Ln1ZRlMHKxWlxsyTWSNSWhUXXNJcux
QusIQiKpGqh+u6gCky7rT1gRnBPzsx5W0siXXMYif0BRotakKDWT0M3cpiCLT2j62yDCvK++vovl
MeNQxjxQokbAYp0dMvNpxf/q38ToJwLPWKyovOLqH2gEet6bibg+lPrRHssJUCZsPxIE1IeViTjQ
FQ1GVYGFu++MvTrqEo1PEErOqtqS5/vstTpsx3KHh14cwikFrvwBHUgwM4Ya6kPtA/vta7B888YR
2FczUHZcQs5++Ya7fXtbeghyqHDwo8CrxLYi9YlRu0st2VGNjCvjUuDWSdB7xBLzv3zc2uWxkfoK
0l9yhVTFmfOJHIkfFjufCXWu/q2dFbXO62uj4M7GTLNHM+BczSt/Ex6v2WIuTak/GNAPMRpLkz/c
9lm9uXaBA4TSQtGCGJlSLz60kCEYmgPMf5ecCrYXFVNgD0yh1dnjhXBW/CDlhqmZ7e0+aNmhw7CB
eFDPYD/6zHSsQdk6yE/g2UoE4pxOdx64ZgNL/TP7I3OW0yA+XRDf8eG9V61vELiSJlIPbJpu8p9x
t5P7fRSyA5RvWwLN0Gr9phrW1X1UIsks9hNcCPzWkaS48UPl6wZzS+xTbezXhe55wA6++Yl2+yq4
FZjs4d+yXU6r6dFWAYb0GxwYUM3wdW/QMNAxS21YsRXTAi4d90U4j0Rx7IcJVvAt1pLpSeO5m3FA
Me9ByguPipiNLqNr9STdKSswPLe5BUm82+gVjqWbr7TnNE7OPLsHFHPXRo9YEfVmjCAoYgnpUOHC
B5B5VsIMxAUKGUy7FbKSkOWjH/aYPVxbB/qznyJWIuRNtl7tm3IpFvKTdyitUTqJozv0D1chJKaG
vHfcmBbSR/DLbrHcdqasgKB3ZDYNuiKMefha+yTlxBmc7mycs6ghPQ95GljhougeykjwJZpHa3EM
Vz6Ar6XepSQ40g+72eFQXYky5gw1KaqO11Nj2X+XvhQ4jiRBKEwb5RPa3nZ1yEDO/Nbrr+DPS1ey
atLujBCMnCEN8K2Mbb71xOdOCadLr2XdKzTExPsl6GwpH8eKYtB1Fi+Uj9px1cByP/pYDqvigRzT
PCRuGENWT+vvkXiVqeiRoa6qEiLb9l9C9FiKuKmiaJdECVv9V0Zw5LqSbro3Rw2lOa8dOUCEwtJI
qPJR6le1dGYEJaOZbM2vKUk02Q5lp72bdEZyLdoBP53hiBSfyHN9SOHytXfxVyFpZkvLdSn9MObQ
2PRV1nofUe2EOKQWSjwAotg2nRXL64cfvQ0kXB8nEfljVYjwGcTrK/aEvApR52zXdgPcVT754qB0
njS13r3yjvSJHJO+O7PacKorVmrxTGr7W8EdGcVFO3fjPTzYQK0aDcmcham1/mhJ0H2hAdnUb1Ep
lZS+szKg+gpdugWFGiNaAqjyEMgZs+uOkcevpI6rtlGC9YM+fb8sBO6mes0HaUtTiO+qrfiaHrdO
ONWoa6DKC5WRPUBTmh6QYyQny4d3sgmA9+klGccsg7SSQPE+j613Plj6081vSe1AOdhfjm+SuK3i
44wSO4zORDPGtV+C85h0CJe5zAFxBR8a+EVZqtE6oHT1Vt/05pYHaLcooedbsvjQymUgj1igQ25L
P5+hfBLJiWwcsyLiJzh/nzz/6SU2if2H5L9TOxz2yafzL//TY8Ld644a5NKYpvvO9I1TzTgr6n0p
XUXFNOmnu0NzC7sveZSFRDRRWy0N9aOmutPOYiA8SluCEAwME69bpeOaIxXC9lJR/c61OYa4YPTm
9Xkc+s+8iERLVUYGBV80LxlrOLi50+KGNFD6obpvuq/CWI5VHjQOG/W2RXSyB/jptwMhWFAAkb5Q
0uBy7Xud5eAWYgOnTst/xYnyal6JsCiOcFsbBnTcR/aXb5KvuL8dOLXiYCUTnldo60f20Z3+CbDg
j5+4elZqoq8EkS12RxLErZXZZpYGtxI0eBOY7IRVcNnCG+PsUO/v/Ic04vrlj1FGRKvhhCPfTsOV
yHO52lx5IdiLJ251UdiwT/gwbmlSsEx/DTQgMiQJxqWpmMVAS3v3IFNNc1wSJdQEvXcCxW2lz+5u
TxxEub/mMxgMojmCwX17TfLPPlEFxZgKzHn5qkwxpwTfI3DPHKrMtFf8N7RNj+Lb4nET/L7s5EzM
4vxIqBqaZX/HUnn6uTkyjKCdvilp2kSI/Iqgg02Bv6REGLT4kHmWdOBfjW1orTT+82E/wINiH0Lc
nx0ZTA7ZTQ4OStqc8U0Bwo8z0YWl9GDVwYgLb+FC5ykYhACuB6M7oepWB7IxQW3cIsjCIASsDlRT
CiGNQ6PQmTJtqzJUVp72+s1lCvUysQ8ODEhBb9E5TI+KbEQKZ6K/AIoJa2Qqp9SdLZh9GZDcztxv
FulKWnjQVGTohjevDu6ICIUQFVzWdHBjPD0/0hCGzSSgt3e4/NzY7wRtpnUNyhkdEdw159o/69Nk
wpCLdgkpgUT05pLXwQ9i9B2hsK8CpDwjnO7flyHL95MfXTr2sIvSGRKS/I0KtievJNfZWEn0+KO5
cqTBkGk1KIpc6dp9OXaLjdm5ocdBuo97FWTG/Dlus5f8rMK06R6Gu3W7m6sCC7Ig/ZnFg+Bt9pGn
Jn6MOChYhsnhT4rg9BOEGM+UYmwWzZd55GbKfdRgjAcYqJUXs+o4vSCxqj3em7OllA/ncYiM8hRX
dIcreAdjMJUOk7S1CZVVTj792JqKEwwCo5jBoGC7DW4Z9sW1F8hcnbccK8kwETo0s2XR/EAP22L1
O3gSDsog5BX58yBXrtW/aepItIbarI/LaWRKedBv0PH42zJcUqgNgYbZGeiiTvcKHj/lgi9QgXnD
+Ud8AI/lbBmK+zbWQCIi8u7GCtL0yMNqiOTA6JtM5gbUBXbrXqZozqRm5x7CW/IhICaANSmOuC0v
zDpW8T2RLp1OyPBHHGfwZjRpV8f3qH62RlCLQ1sbmbwKG/NIdKO5j+tBCnTZy1vXkpcNJ89po5is
YBjFozUcH3tvbEeiygZ9YGn4Y/a9DsuYxLrnBUcv7aQgmsaFDQyyTBdaCzhUUbsy1OODBaNZx1+E
sBSCLM7OaKGFTFmhVxiey8nRQHwomZkZy0jrzoGyRFkZPM3kX/lYCge3xXbFlOXf0WBiYTGfxAU/
svBFn7PBvNrlFBYP/l+fhpxO1/xVMcTYzUD5kPIOQm+I6qqUexgdATM4x9o8IOYPSCCv9ZC/HOzz
j6X8AlzeFsIKqTMuFtkvJ8f5wLDDRLqoXpC6i69bOB+hyw5rZzB70AtSTPd+Gy9WBAcLuEO70sNh
FrrklcX2YtDpz6JWeYA3pkX3b1kLAtfbvtc4aLs/5X9u+Z5TKmGKWwFxBeAF6auQYuv2Fa0PGO0y
h7P1tdFfzsr8B30eR8sHAoraPIc7ypyxM7CBVvEKHw+Lz7ct9CmoR1ugdUQ2rISDsw2Kv4wVInGm
5xAmIpQDXLDMqL6XksqeMb4jmvBwevRDSXm9KJW5E4IW0i8RHYIPpVRDb5qwVWN7k3ak+Vz5m0vX
V04NXnPBII32NyuPjq8cDd2xPaBRonjLrNTO5goaVbCSai68gWkbikkKUxlc63v8O0hyzsF9Swpi
mJF8hTjGl3L9Vm3M75W0cDMLwCEB8H0KLATmeAeRlSd4SNZ22bBj0+8Z3MzLnHCpp8fDbexZQDKS
TBKyGptLCentq6ScSAvKXhnIaODK8V5fJODWeK4G5fpzToAJddj18UhOIb3XP55pFd9KFqArnIPE
SgL69lW+GAkAFgqe7jjcfkPJKDiywZr1W59SIEfddTcQ1VW1qD7UR4RJsM5Dwq76UR6FNfR5QVk0
OLvJq1wQLvV/DEOPNL8nZE6v9oQRpPSLeKfACU1TUGOBfiK5ofB86YPeH4KYv6uDZHkptrdfQK/J
8CKGIy1PHHkeXWIUwcigX6ySUWTCido5W9K1uUyE4xJV4+QCj0trlZz1gtdOe/oEo/IFeyEtTNqa
Y2okdpII7+eMzZDEvNSVPROmmeXToKbizdig+gEmfocYSISUdZLYgr5TiTCb9FstbdIAfLMygXRq
9dN+MbhPPJIFf0Tqoma/gpWpL5VhZ4LhBmUm2mLNVu+DkbzvWyc/7WclEfOPWoYiO1Q1HHjVgua7
KXWG5NYmC0KG1srZmyDBbsZ+TB4useA2pB21Lo/4IzGLFXFsI5WtPToW7bMFPrEqd1mhYnDOI7um
B+WhYxdSPRbfw02FdyyPZ9s8K62azoLUpLU23tz8qzszjS/X1FF7dKEwyX/VQ2TztWiHeTXBY2TW
PyIApFPPAVUHYycvAwvuoiUHv/qdHuRpBb7nGZ5HLK60UNOLS3X7BWU36E83ziq3LnRSJGu1qvKB
pcXzXBSjpabc6WAMrricAiEpWJN+6333ouApifWSsBWCrd8BT94dIj1hIDYxvcjW+RjqVZhXBOGR
qWetFn/SZhvdyKfHLmyEYbv6nzMVlzYLdN3+OGvwZpFCYOLGPxVzNoQI3MlASs3MIbqU8fV9y1he
AIyvG72oerGVYyN70CAaS9ppNndQQpkLq88huGk5XHnReo7lWzYIwFc7uF3P0WmtSqzxg/MxU67E
0ejT5B7nBT4Pig8pDhDJrT+ldd+b4DRsRQanrgrauf3eVKjFaD1ZNIt6Y02MfbOoam41qLvyO/t4
Sg36F1SHddNh5NZakxCHEe+CX5L1w3B155WSFYFdYkchMuqi2KIjUPPGxiyedbOygtWtlmHnNR69
cOcnI7vvQw6eXRCEVlVOhd3b524JezfmuHa8lo1g9S/vFXo4L4j8GgTbFSeavl3jAXhrAj7dhhRx
Esxm6KAufakbwCChZiJA/nT8x3dCM2mbzCzU66V6hqzuJcQ5LdPNpvurvYHXeBwLILVNK4k9a7+9
nnNxY6eighqvHleeFvIuItBl5wpeHjDiUDGeJWLSfVwXLO8qWimU8S6tXsWZ6FzP768U3TDCLeTU
87ap55Z5BrQzB6UX8aJ+5I+4qMoJHdJN3L5LZvbHyjUPcZhXmYEKguNeKalna5H4cTy9qS6rGyvA
Qc6qPbCNdnD0LnVMVqDKO6usR9njfqIpeTbokhEoFKmxzwTdNO8WL+Pz3gbz2VThkv+ozC3oWtnx
XoCr/S9UHy4p9zI5ksegZwLOGpf4tDTc5wh1m5/B4tGNppJTCREuOQYpiZI8rrCZQE6e/dM8SbQu
EOTMi3x+6kR0nkLlIEgmGVj6Uijq9dxoCodHpusCL3nsFfsC1vGKWfV6mtFVl44SSDXhlSc1AKc9
86n6pxKcj8ZPgvpVWp5jr+46DFjoET+y/W1aczsFeLuHXomQWni2MJwbW8hmug9e2xDEzq4juIxI
QM1Iqb3Ky55XtuahcFqm40/GSwSFqAkgpzN78wLH6fFCxH+Lp4tEuhtdtmwq50lNh5ltq1/O3SzT
ASAjInM2fvkBZ6IVh6eP3h2KZNpudhzfLAL8DNe5P59WAj/8QT0cHX8rbFnyWR2P6gC3N62RMys2
t4cQK7mjD122wHI/1yYmOHMXmzZatBt5VN+Flc+oBcP0ZyMuxP+Js36Jj29c7vZ8B496/CwktrTf
MoVVCkc0s8tYgUIPQjuLVuNiKa76NLuX/tH99gAoP2ZCaPK750CVUqCA5ZIgSX03d8S7ZyKjhLj6
0ZmxlRLJ8UUm1pU+71KvRr980qSzpLVRXfSX7wxWYgmO1LArRGLO5ED9qHWtLeAHw4vROeLzVSpU
Lxasah3sss7fGadfLfC9dMcF+lvHBz/fmbufw0bFOFilHptaHzrsbk6k4oHs/ebVbfpDm8mAgHPe
b3eQM0TJizM2778S2NA+alqfAEpiR97Vys8DAlrv6yeyossuSPmfO1E+52EXfpZpErXj8iOSHhJD
Tvzz1dU4HP3xe3Q5E3nfUTM4CvltEp5qELrvR37SP/g7pMVcRSzQm3blSeS1kdauYikhEWshNHxy
Ay7Ws7wkQWc0PXWAzNpmKZ8buKIMzcCr4RAd8pU/YheSf+iynuQhbOdhJIgot9kzPWGXN4dcJ3W/
caLk82UG7tNwWBCt5pD3h8PPgN6jh37JUxspnLdi7vxVRDHGUZpCSXWdyyy+NrAxH0hHWGf7HUn3
pW1n/T10yTWyyO468MVdGYViuqSRUIgIm6tf6dXNF7fKcEhRppklIsycU3fdtGUcmOd6fUGZZoLf
2VW5D2RI5zo5qYwCs2aqYAhfRuGM5/9nBKKfwzx2Duig3pfE+oplKV2c1QTAZ+aV1K+aPUSis0mj
qa8ss8GlRfQkHnC+4THR8tCfH7RA/XcqVS1dsnkxGMVVIKCNP/pU9XUv+pFV6b6le0rZYOmQ0P3j
vtFwSQJJe6fbhjE7nVoFrFM1E51q80Q9V5xcIqQho31mYw4Dk+2nBAFKWsIHCXHAKFHodIdjcBiA
PX7/yCp+CESNInDItO7M+uhyq4tHQvC544iKmLkQEZCtqhPPtdtV3lcjIM6tyM1XxaGB/ZKbf104
WulzDXYwUt9pSkD3jVNIydBMX0X1z3gQLP4Ju/9CzIKEexr6fwLIe400A5/HTPRDReEkuP+RcRF5
1Un7DVqbtj+L/MQcMOyYF/DtbE6nFTIXHOJNe49KCS6pCR+IGUGB38jWB6VZhXdUt67yWu23VgMA
8857+/1QFWWtDKnaqenlhHHDqUcbD1eWq4sg8aLgvY5Z5jsSqeykM0EmEC/aYjspwz/d7aUT5Di5
Xxgl7gis2pvLzDqnebul3F8mIagKOHlmD/uvvFygFMLAevgYQO7BVkpIRSyJtgTR1YA73Wgqfh5H
TmeOjenqCLFOnCHWDnHm5TTuUfy5H4jZcK7oUM6fokRfDWwmCgkUG6oFnWV4qKpQL47dpZ9EwryM
MS8j+bE7WtWgIN3C8KQqkemCnR8ze5XIPz4vMITx7i3PpknvgKxem0XFqz1rXFZTfL+/Pev6O+Mr
CwtvTiCg5mIQQyjR89UZEgR/HRwzfjFXunzY3oz9WinkfTbLDjxtvbU4iYGBIxoDv2LHlXmlJiV9
w4ZOv1Fxp0jGf9P1U5mOq00UirBCiHmHbdY47t6s21BBMgOqJOwBb8tDDfP/doSUgN8Ai8cLGkXT
0W/7g6HDU9nmUV+8T0lKhOW2BgHYi5g0LVa2dhQbn5rAWorPXFlrQ/1rHFxm8mfEbgks7TcQfJQH
icZFbcI+0phlCv2/zzeES1fUeo9hpqU8Afz9/V2bPOnwgM8PisO1pGeJ0MssPkTKE9B/ujz8OUBM
A8Q5BR0ulYbiQ1sgWEDv7BVJtTa93veIjaq2JG38lmvXbLx3fyia8I3NOS+SapQs/PIC7mKu2sef
Nj1TYx1Ui/gY3VRWZ3zu0lMR65Wwk1zhrxT1qXmBzL1nJhxqO0QDcvyNjGyXrQQ374U0hdpPVktT
PEQTTqXyNyQ+OP7bOVYDMfIACT/hNq1uuJU13Ru6N/hxMNs0yf4/zzrvSnmXujrhbC67sEuVArtj
+cYLnRrcP2Z5ub2f6VPLEcUuLZJjuckWYRDf6aJ7O8vTZ2p1+qN07Tt0JYmf8n8V+HxXQZIhcTtA
mqTLPux6Aojesz4ZkZFw6qKERLekfDgdDGv48cpRCfeHQyFSJ27PK9yChJKwv38kSUsGvU7OOf75
i61U/wOA0RXltcgYkqZ18Njd5xMHTiXachGhL2h4riarnhg3ybtu3LlBsCMNRpdqnGAPtfxobN6H
AkphBLc0r9e6qz396M7q4k59bqY/QtiAtQXEah5WW980yYuA/MItvjsOi00LjmFtV61NQrn202Ki
geBDl6Bcl9fZRXeAkgjvmfljyKzrsrPDxr4jtPjIvWrGyc0dvSI8xiwJLA3X4cfw4N/lr+ResKBN
yj/DZhyHLA8H0kv3JLjfvtVm7pDWrsdfUNzyJfaIuw5wP+DY9jDOTxleV66k6SXZlzHvinTnH44J
ZKYVgayjsxJaT2DSFZfNSV8MsQkgecsS19np7ADwSsn1B/UVlyI+TRjECW9S/ZT3zD2aWuHjtU3d
vbgDMVWfFlZbzkjATKHl0CW0pokD9rTPYhb/VwWIkXmb53qWTRJAegdLpHBp3v42Jh16eVSWvVaD
cpQfOIczS9jOAE2a4UvsUdIxLWn+ITj6IAz9sXtg97hOG4Jph8sFoYz4/0mZuL0z+U8yvnNUkUof
R7eZY1X43trW0HvchSb9RBSRuWX2NESgvqy0phP32pjSjM+rJQWwq0OyHJtONqhMZ/Et7Cs+ftMt
ZX4j6XymO52nSIAUNnDzFT/iRbxU86zOOKBvgO/BtJ+ygVRO2rMpPkcK5qIOk9Q0f419htg6S9Ku
LF89JLsQ6wDjz7y3TsbGtu0V0m9t6vgSryWgQYblhXOmgrMgxvn/5EEpU2g2KLVv4k6Vr+3+Soob
sMHJsP0/7qEZyx7/BmhOiJH9GFmLAjx36pomYPCAl+QOcu0hamnpwnJoC/rxMkiP+0UtHtiikaoF
RXSm5cDHct/A/k8+Te8VmXVrIUj2xLBnyFZQbMaOt1XLMRzQ3ZsLcdAde2nz6V1OUwZ7YXluEujG
IqBxzjgQawoohuuiZ+EkMTlMqZgTtTQUPWaCKFjMRX+VMKQfKm+Mdrkely//OlKp2JGI5opVhQ14
DxzAmtJb+O4J6T7xyw4ALIunydgCQG1gVxTnXLgOqoc9lMWVRZs1xZTb7xgHJGvLrRthNwICsqxw
Q/JrXSw6ed+ptGrT3kMgH3rAsjVLNFSmCFIFAQfrZz/Ly5ZBLRis17yFtYw6xWvD1XBstX/SiW6j
kdIo9l3/2jl6hNZRiwf9DXwbCFFkOi53vDFr+GRkrQw3LEZcXNzBqWtsIwlAch73ejtnpRXvlwkq
FCMNlnVvh/V/c5XdmYWivRW2XNbKI5poJsaeuKr1HL661yDUeglPI5xk/e+8VqhkER3NkyIplaTH
E21BP0CRTwT6xce+6ky62htwndT8VpVh6hQuEs/3virAAVEH+2SmPve0DlTJ1KOjC1qGClI9P4Ay
tiH2GwwrGcxsK5txGqGLgnvXkQ7JocL1RClLeHb1SVmoGKNS/hmd4O2/BjqfoYNz8e8jlvBYqiZO
pG3rie2kkXfjuK43xJ3wUleokXavTcqLPJk5z2iFn97TgB0cr5KzePYwSeVtxfIGEmBs7nHiUAKh
pc3hPhZzHkR6YJGTXW0rZMgtfn7Kim0Xlk79gfujJexMcdmaCKAj71lSqGt+uvDCeeUSxPv+7tUK
pMW7qkOR57GUOuVVk5ZL1iSLiMZehA8rstua7VVE70s4RPhyQ8ibumkyzDeNaBWdiP4uuyW5gkjq
l+O7qzNlJT4+mmXetPo/VIdp47VmX45xqDmsn2CLnmXkpDVk1yv9+bTZqGfM8xlNT+wwm8KuWgGT
VB1OfCPDOnNxX3x7F0cd/HnbdWHyWn7zgvkkSPMiWyDo+rPS4tFlmGZEkZnZaRC3L3c7v33kBuVT
rQGeC9r3U5VsdcY5q3BigMIUTgjoVmhj5qwF8m1T+jL7+kUZDNXePwWr1ri9OJ/RG9oMk8CmA6nL
XdJ3p1gW01iEeRFlIdZeuO81Qo/uXh8X0SXKp4CRulzlvQSRI99og+sBR9QP2XeoNSM55vbEvWfM
daPTJoNj+mT0oE/S7cunX+J6+oDLUwTmC/uivcqt4ZoTFFX9BSeSNqqW7nZ9FzIBpNJu7H2omxHh
07U5aSF3QBH/b++KU6gPwGpVI8K2A0el1J2dLQXqYsvAqz2Bgq52PsPc0UpwDEfyRNnTqaJ/IGih
WLL2ZRbbmL9sWxuVzdvHhp3zv310QC8W4J/SqZIM9RKSYCRAK290FzVaifEmOSfEqkh8eZ19RktU
C+XtOXrYs5dGoOSUySqqtmPIn4QVfIKnJ+E7Wd3c2uVW+xBGGm8KbGJhyVAiavqivzqTcLL7SvFT
9TDYfv5mZThOz03P1cw5S1C5SSRNTu/6cBv8O6J18Rfyhsc6F1Nz2SSoMZi4S7bU61GYANEJCgMK
e6NH7J9A7/Hl2hRPZIBeWOJZOU81uhIrdYCVpf0Sw2gqdloYb3jAE+h/ZMo+Zz3FKVnK4YYHRx5U
/LWCx1lzH0Q6KeI9RT4LcouZggRz5WTdOrlz+k7Ht1ev5+wQ+pO0Fl6agJzozXeygnrHHdQFxklX
rJ43cjQ1HVL44499gEteE2JzcuHlU5X5UmuJFObh+jNnAtc1urA3fusS+b4E5N5p0AEW0lHm5TGx
LjdimTRcA81khxxDMmfOVvE/U1RMEbet6aOol3qWo+xP0UYzm19O+mBGGw5HaKDzYQPjboKMhccx
F+79vruCBAxlKgNe7F4nyMK/Vdwy0oTveGahQuz0sUubtRWF9XtVz2lXQZf12T9rcPUbCXfluRx/
dR0meIB2acVvTSSSPU78dhxI8HQW1vVpx8ymReroeT7sPjGvDKbzbsPwAtNrbKyqhjf1KIkpnWVG
OQkR3rjg4C/ekEgTBu28XDBoDkyowjJB5OHyNfVPp1azQ6X3IaBKnIpzEYIO6yRc5JewiXy0p4i4
0rtWTwjeihR1LvdbK8u3pX0aZNq3z2Ikxwne8P5g3ayKtaeXRG7r1jpmANvCWMJ9NXzxKgVKhkJw
Fx/IiABXzvn8P1llFRDF52PwQ78avRx2OosrJxpVywa9k8ZUly4+YV7600k+xZAOr8b/HL3K55Mv
gBJUS2Hblc6H0j1J7bAR4MtlsZGO2isE5gsFJqd0rSLTl18KLNe9IYLA0YnSvu/tLI5z3PEeV4RV
lMLnIKlzaXT4xbi8ZBVkaqb0WpXDlUENpKZ7eNOrn2i9o4D5sLYIGYUIz6LplGsKhxVNZPmyKQHX
uwBkHy5YxiNGmB+NBt6g5XhO9DwW7BdhYTPsMFmtdFrf1YYbiNCsq+728lFhPFaBj4d9eamKloZp
AUXozw9UL+uC+rC4dbe6mZim9g+huMlu0jX9Ba07YcIoYmKgXyTQRCQ5mX+2Mz4Ldu1I1qLfeNX7
8t/JnbL3zpnoFAYpXG+PAzIwtk6IyKb2xzwtV9vne8JGS8sP6tukvw9iaIjZDW1tgoWx+Js4+MhO
CNzlRFoVBBozrcAQyNejR9cjkHBK07TnTOWzhiBnZvKARkN72PYz+T8JFgIk7b+P3gFGnfdmr6P/
0odtHw8Vmimi9jobxUYoPIOLdtmgKe4t6PicjjGkqCXPssTwSLGNAHpwhFFziXxiQzulzKekBDKc
yRcBGKpRBtWqdvzPnluc5i67wvEzrn4Rhz+Hx8navYS0PYxqdmLqaYZiCOsgnQDgbUkvGXNTNr1i
GuYqVQongasxiWMWM28AssAU7QMov3qVbF3sAG7yeQsY4mj0hVbM+lGsAu4EIdWdzrXA7SlxkdHJ
ZI54lRhlfKaswHS4L/gt6U/CUEJieoudre8XRKbVUbqYCvOCXE17EnZUGUD5HwAEapshLGW5yaN3
JF6DwGxKm0BDmqkxQAmU2LWpC0d4VcGI7Kv94Hfg8+uJnsaQPI5I/XOukWHt5uQXfzKsAzruSMOz
ynFnnlT8LolanM2pX0WTgNDNnUoPAm3pDsvx0ucMjBKqPMxHrSEozuFnjk7TBsCPyHQbOoHGd0O3
S1XGruEtmWxRspz87kyg0KSYAwbqju9tziaoPK3Y9ExAtXVWAX0bGwQcupnTnkq1p6OTPoRoi/Hf
mNwh8nzaIIIfaGatIgFd+e0avTGRh9jU2/pi1Uz178MU+fo5ky70pJtQY7nHgeW7akevxNbXjBrd
moBaR08TKtLe81bmv3H+3RD150RZSzPXdC7lKB9OZ6lnnMzMoSY6DLInwg0br6RtqSm2aS4BDMhK
NCKURg7H8yvChPxIC4iu0CCqvFWdraE+fU15Jr5RUk/erRi6R3zslZyRC9V9to8TSSZ+ehbTenVj
G4vS09xlXUE8biP8KYKBfSnxmEg7DzwIorYAjLs733IO6Ii7HE1I+TQZYh4MpqsaA41W90u7STao
qRN95B9oTEHwdyi4+qaTrSYJypBwnk3fzfSSCd8+G3qS6zrZ5QrNv1Hi84cNAxIT3XQDZ7YHqzgi
bjtWyxTvON6tEyfaRuQjHxTLKFflv9m7T+w1TsUJ+T/TbT3/pB7Zy3Bd2y3ayrvnNqQ6ZZhwKHdA
VRkAfJanfXDIlIarggKocQC7f9Vs5dIkEj7aWbzSINLdF3pm9E1rtdwlnBFq0g7+e2xvy1Cbww7k
ZaHrJt23L1g5WravxMfoacoFeDWB+3xyliak8ktbK/yEcCBnPcyau7LhOeKhw8iLv+mOWsU/4gvI
7l4tWnDpg9015wEPOnZ9PNqpdi/1bInM9oZoMa63cjex4ZWz5T0e8cOFxX7hIJXL2SegY0jls65A
4PaU7vjsyLcaBYHz3M62wzv/eVKjWMML6TB8tvdHzQkIk3nv0KrodywLWTlt+9oC5ptT7cjwL0Ya
3knDVPeiqSVFojCZbBU419gmaNeYzx86tUnwnSXjg9fKiMuGKeoL7ptFwxvGtkFO9buM3YLzKgGS
10FisOpiuUn0748Ftt2o9jHhQ80WN6MyVOu4TsO5dYeByQhKfil4V3U0rW4YzVtew3ZeN+NYfvXc
LO352062uoJCJv0HFrntxLdESvWyaGwjlm2y+DLiGXGHsxixFDwIIJAGn176sXKWHePz4Bq+6xzH
oAzwsmnxnkT9/Fa4M6uHU9Pt/ijC80oCb/ZQt6YPDIElQxRZqdlAtZzeAaElBOdA0sY4kqtDgCzL
rTjyYxNosZDuLr3OqfY2re0ul2dYYz2v8m3M9JrRNEwoveaP5MqRnL3E1xD9kTKYFO0ZMlfUy6nz
7le/yvv3rov3P8wnuRT5JhDAu58A4t6mAwtPTNzI9GvhUG+pIH6vcscIG6rQTaiaMxevcIrU3ke4
7yWm1U/1mzVhICjM/cSIvjsYB4AH4OeP4Cb/6wqHVQr/zCxAYWQCTVirljql09dCBMjEcLVG9yAi
vM1V9LLlBWqerZOXX1lx/p7pFpTXyGH1My4Mwu+yc/H+tg/uaXOYJwlVL8mbqqtW8mkeUngASATY
PvVVTfXX1sLVEpYbxbysPJ4q+aPNLkIVX/iVY+yOA9AVO25FJXBAy1/Ai1JRDenLVOQFSYzzC6g8
24LOnu73TPWfrO6Wju29M68zeZjH8vltzwjY2jPmWbV1Qh1yW4hfdGGeBKIcAtPaXOSRHhNr1YLq
EBS1SNmycwKvGbMir/oL+6+JuPH5gFrTdmwnQgh+RWioIA1BelJUSnXJ8/ivQrwEvoisyQSDVz10
es9UkBZgamxH+BpUUWmEAfJwKlX7sAN1X58tue2gneGudHkcVasQlKp0h/oueEhRuWVeCEeJ0LnW
PlyqtJuPLsQodLWecVzEY8nHTeCvGoc/Fws0PxspNMoAuiwAm2uo50ZLCrw3tUBcAJiSQJnM+e5E
3APDhCwvl9GxXohBRkvmUbiUsKZh3v1/jJN/nmeaPux9WATuU9yLjHP/JMNdvlUa9Rdh3Fud00t7
ptL+51t8SetN7OUl9l7EOD1nvw8TrO0ldXIgjd0zFSnZwgq/bW5s+gXd00IZK+WGYH4H8gc+NrEW
sTihKSUWYB4SAohM60pifJVL4AwDYRZWTvn46Beqc9He4FCsC8HAttoKUIosFf1hvcjnBDNi5kcd
j5bP3H+crZsvInwUsrEYRXR4npSBgAmgsdg8l7k+3lMuXSg7hC6LlMhic4XNlHjapi/YgcJwbDCY
Vr+x2o0RKk6lU2dT5Pn73tgejZDhHKH8rj74ASTeinSebIjGZbhPSxSgTCqd01sPD12xf4awgVFN
kHUE5HZkuMHImaBGfkeYA4UCFClRPgyjtbV3/TTfBcFwGiI8ZBhaVzX5wGhzX6jShBjFb32anpM8
yzxfyWn/Enlu6HMUdXB5n61ICtw/yFbrDD40iJBFiAcJRj2hkGhBdf0nmkzdYmpTE1NtqpbYlm8l
CQKLSVsgY1rj/f08QDulXcVX1f+BAgNBv88z/iQVhbTOlH1eusC49cpbBPosE3NUgIy4KWtG7Tl6
wvLo6OB+xAtlIPHvdu92jNKPwwmhktOPvsJJtXsaQcHQEYWxfbmyzjWNsMhWbtaD7hQ4x7fNU3wO
/II7RKp8Pd40cf/ouUkkesOkxAG6vNtyHb5QQM8/bSirlhU+1KH+GteK5hWcsznop5idbgLrknHL
Sl+62iIO7XDWtQXNDrPZMlFyYaAN3SY7FV5VOKEfKbn9OzqczNYzbSX4uE9DzgYq1mOV7t3HuDGT
hhdKdJr8oZVKIUilYJt1pivbA6mBUiV9vpZzXeDjKb7u9S6FexIM+OhryTsSmIERHR/ZnOyBw/Pl
yWLEpt8EXBYWSbrOw511lUayrZ+jrIVsAF5eFGUcXMn2UoV8ILr48iAq55ZlEXRNimxy2SP6FoG5
dBDv8/ls3ygFl8NGgW5xcLo/CujzE7gz/FBm+0GDjc7dt28fln47YP2l+LivoVIlMHgOK7C/b5YR
4YdWmpXyou3A1ld9d5nXcVzlvzjf4c8jthEfU7IkK9bU9/zxco445aJh6NVjJ9HIjry3RI06LpGg
VlE2PvQWKJ3pWkekXMRVpgYdWkVfZx2k+D9lLFp+wlhHYVUkGbAIMJ8n3Q3vY/sFrPjFurT5nTIm
BLw0j/BKqKsMTogQhx+WV/906Ubfi9GZ9DcNed25vg2ZHX+UPfCIA42uzY/KLCg+ob6mo9lGIjba
fpmkoTCJtxjtMiUlvN4730WZfORVwFWPZV7yDcVyAaxZN7fh8An60TpnmUrlruiHYuIY7Qwn4+pY
uo+OJdGg7RBvh8KAqVp0EnYYbU6kBlmUbfLCu/MsP3+koLIzQlG2XOSs2kqR14fjpTh+I8VPeKfJ
bwr6Q9uUmrxbjj0qMxklcCRWUaYvJ7Aq9tRy1jqzF14wLfjhClhld0pfrpHF4oZTOKj8TgysUtxz
mcYVaYXnZJkAz/ONL73sKuArWqMCnHiSwkXQWt9zjL0Zd4Yam3JAfr/3A9ylYkSwSDV1p/AF7jaw
BOQnEwuaRa4YB1TA68IQLsdbZBJtTo55e/40Zc69rIwyHWeEdM36vgbVURGmW8Ba3Gw02tEBt1yq
eWvfQt2HBL9pZb4pdLDwQu4qe1BtjQqn1aw3AMEWcqu7j9gJeF0QLJPrmEZz0GtFbIkeZy4Dw8vM
/Dhr9DOh6C1c+xGlVnp9Ov2XzmrEwaTpZ0NeJwb+TOtLTYUkS9cVj7JDqIYu4Wtx/wbGSiSgGHwQ
83BJ25e0ZEyep2Ex8r7GmMZUvzguaih7NbixmMDLkcaLj5RhOf2W97Bw4ZKmOOPn40EULSmzoSpZ
WN1Up8yAe2Sqm9dJKsVbagZNZfBeCiRitchHSMbuykXyu32cPWMOpPTw4SaLXa2fPYzZ++3NW6bO
ejEf3tnQ1RPQzgDs1osMVj3cj7pwP8GQmXBeb+M26Ioualm3O1aZlQPguzxGN8jLW6LIaDtXMnnp
xkEjBXAg76ulcCy63UXWLHhD+FWgIu2wtmKVt4JHbCYVjhMNpAdFHxxj0Mm9XFW59o7KcpWO4n2U
L6hls7tmdr5+mrRc8/OV4gBEPq3awWNklRFY+myTMM3/hNCcFrR850rS2JvVehaeIjPwnJhU7L02
POBt3887gAqt+MlWaBt1Pl8Ft31yPsxQxcgTQ12s6dBsBaLXVYYKKHZLrGlsO+19hREFuodckaQ2
ZGtJR9zeLiiOl2zIHnevoiVdQAULhQrp1YKr91F2eiidPEtFkxLktydRskePKeTsCPRHoYL2EM6p
RXAIpcdGO/ts3jkQyWQa7fdo4XgsEQz3JOUn2AEKem+ESfBzgVGJ8jcb1AKVKY8xjzEqMoeQz1Jh
8dfxl8wZ3PMUc9NmYBvCuFxcxIq3hl/GGQfAf0H69+kMtqE0+sHfQMyby8s/RJWE/4ltVA2MVkRI
MY2xv7ROhgj4EsGSmC+n0QofsBxs4d23F5dt81ijZb3YSCxKAqIuLfpMmpipEsYtGCGB4f6R14yp
K8zjratULuzqXoB0F34PLMJZThnsyiHlMtz/gOMbE0FTuUiRQa302Zh7LhTHKlbi6dEa3nVA5ZzO
yb9IMXc8s/FMcqJSfcJOqFq0JrguXivSMg8gvjgDOPB86QM/41/OXHuFKgVf7AeCmtHtkoiduP4r
JL+TPXLXyhkC1OcyYRm58/rb3c9sKnJQkMWceRqA+yll4ZXq1zb9UfQbRMcT78sbB4ufOTmcm7Ki
/H+tebpvZIdCYz2QxIayd+o0Lxt7vjRZrSHrigSAM4omSezzLiAfZfHkuXOGu/aqzrTK5N8yJkBI
CEQUGD1530zzLdq6PeQsFE5583T0QRlrFVp6B9RAbkMExu7035qPOdgRXafa7HcRaoNXtjnKtvPs
xeJzNuLGyybjrh+B5kYc3QMuv/Kp+jrfgq9dC+SsqenhXdLURRIt7ZI6jDb7IvcKVDW8FpayJKp9
TbNoxYRc2S8AUBp13AZXENbz2p1OeGQXe6UMvOYYEWBbreSQ7n474EmWLfTHKkKGiCv3LTnNXLJH
hBKhZGzmLTufe9f7dU1Nhdc/6DFGZF2QA1mU3i8rZWERuZ4Vuq0Eg+1zPZjNcNjXZqIKDb4hPmtj
0fA3/PfV2d+62KxaPuRZwKNmmtPBv3UyNBnoBr5wfOeHK2D4fjIyBhZaHqtGubPUqIU/2Z5GNDBR
hVbuzzVeIrpKVVSBkIdI9sfjUvsaEfnDocpb46p/wdP9ieu2z1Vx6bWQGuWSHy99fZy0e5z7PH34
IyyQnMLGRgox6BR3WqNr0zCjCJdXzE5rxWbzGuwwYvTWCWDCcDNqCOtIHJSqXirMqSSVG0v710it
0p+N7+5AlAGEf59RIIHRrjrZlmqbi4hZxOpaqJsqBYDiGDX9Xmz1y/qipDSTchFOGRIgrSMpvHXS
QVsqCUapXB5vgFXqF0lu3W6GeDFAlhpFk6kQW3mYJOdKO1JsjPhTnSw1XD2XUox8Pgq9CYbClqKr
rB9vtZJXwfqlKqmte3CMghVs8H7grUbrJ6o9UkvoCf10Ta2C71ofvpCaMM/GcWBPiQlg2Ed3a9IC
rebLZoxJ4wOoXyRVbqmO/KNmoo5DnxIhWTH0wLRgHjyVYaoJ3IKyMhgUjyTefG0QTIJPQPNjG61u
kGRHq9gitSqnbyXTQUB5QyJ54MrEpW5zWpGsWGlTr9bckK9Vk4Cm5/ij/sBgH8B8+1FpMyfubVpb
0tQGz1LofgO9lipWyIY3ucndZRcyai7mBSMmo1xhXDMRuXO+FuPfrGnIYCSKXtrwKe0uBzL3OKBE
jf5rDYdpYggEYzp3q8upEvrbMvnvq8dplwV0R+Bjd2NI7exZez1OdJ3I/Yhaw7IFN21deralb4Ez
hCr51fNVUMB0zV92LU1DpLGqlwYk743cv70BHQ935yD5vBOdHEV37Zts2tyTtZsopairNDjalm4Z
F2uY76EYBvigpTWDrqAxSuIDR9ZTFHEij3aUfvztNTsVifQ/zm3weAn5BsThAPc0Bh98w0pJ3K8o
1t6f0rKkwRJ8g5dwswjGSiYtO4eTMoFEIqSUTGGospV0e8ZRm6Xs1EJJpk/x4iSLa53jH2yLhnhP
YN1Kxnb9skj2BGddGH/H2SGS3QhWckLP0Y9n9d7HpUgWRs2TOvpbpg2KmW+h6b1oUVx7+1wiCxVW
ntq6+0Fci6EzxFcBmDMSgpx6Kob0tHLkg1lVq4dbTQnFnPtNp1c2U4uoBU5wR/uJgC6y41XsC6vz
qYO1I2Bvb3NCJSM0/MS51Mx1T/NmqoDB6L2hoSOAYPFYzQx3dUVp6OEr9mQvUA4w48eNVHtuCy5p
sGNS2heQ+2VRKo4mdk6buTv56moh/Ds5SvwUWf64bqrVZ62nnysB8WLgy4O6r7c4J65PnMiZqFDr
Qdh6wJ0KqN+YqgHk2k+WNYdh412lzbhdPmwP4wJFV/bmSSN32I07+yB3v0hKjiYUReMu8viKHana
EIDt5yjtUWnG6mtkmb8jFmI/4xfFwmP5JD0XYsPOE9JgzM/Iyz6ieVIQSqIMDbUw2jKgeHUeQEfx
quIw580gLXc7VJpXlz2n5H6tPXCXC7MnNG277TxLT4fvQkZL3F85qwXzshldcu3n6SrCBcMGIb3S
m35fYPlYahiOg3EdkdV1K6k53d6lJc55YtWHYLromuj8vHR5NKxSf1Xiud7iw8OpEM4T+ucg53+L
BEWxAgFIbcQGo9vKLk/kXwPdwEkDNVkw8DtFDFRBGSNgF16JLve/7sCFz8vEaAyhGTK7WBWnwgDF
fA8NgF8eRB0ratLEfXJlEMFTl6VSQ3u6Nl4z0ocVKQyRQuGGwRxAbUZO89I4zTMC8b8D65Wa+us8
iy2h2pe3WR7qp4BpWTNKIjnrMme33Y13cbwxZGCGZaAM/oNRsnX+aSAbFpnd/OiA/RNP1E28b64U
2s8EwuhVupqbc2vBhTvHO0eYmQIcTiBcu1S6BEByxrZxUkvCT5L4kDVyT4r4LxBDGL3b01ZbOOLE
TiAsvaH627sH3CWKqqGPjxn4ZpCoGC+/XJC5r0o21rOL/y+44wV9tL4lP077TrspxVSEpZLz8iKo
n5w9r8j/GeUDtpFIzWpxlJjawJZkqQSNxVGjl1iklwdsIB+3YqL96G+gqebFj7h5sEOeiZCBUwzk
N7Uk1Xk2XNoCO8hx8KxsReW9kXezLmtwzQCaTm/7tlO4JKjT5bo3ae/1Ml2wea2k7/rsxKGXA32W
3WwoNyknqveqhooFjEMA2KBrGaFqdBbA5t5cf1/h2m4qAzlLFGAbi6p+mim2nrCK+5/B0OJVS+Sx
eaAb7+Sn5IM1YMTtYrNglmGwWZY0YurEPGfZfyb2rmw5fo7vCEwQm8NZHb+em7DiGXhzRwMOmJZS
wNNMJ+hHJOm7bgfG9aahLqzBS0Qu7/UksmDYjUqJLGiOEnuOlc6/cWjSVWCcnNQl3uVjkOt9LHDt
Db6CSBMdgdiwBanF9zrfqHAjTuiGoHhoCmI2Cr/zzUnosSdA4XkZMylr7n2FoFTAWg33JPTYwF3w
t7+FFvBYVdFicQcCx3cga4manhQM4gPu9ozNFZw2KGe7mVTmiEXYi/8KDxJF69nysNHNAdKUM+cp
7KXBN4w49TFL0+9snx6dBNUXqvuPReatp/rUQd763D3+3tPxszEd9t/Eorujm7CPyXrssATN2pyZ
xqzmc40ioSgw/wjMeH3pcON36tRcill675acxyPo6ErZouNBkoXFj6PUzxZD3j1Ym4A2Zz2ylD9M
bv9UCaQD3bazWfjziXH4KBSrH9twGD1r/3Vu2pGRYIsVJAay5TtCDty6KQyjrC6hMkSyh3QvJJRL
4yeEph8DvzK4jDmBZ62eOxIPQhnYgjipAZ+QRV33PiJ2SWXdBjreXnI0TOcnwxsql3zoVIWqdG8S
OYZHbhHUzgi2Fc032Hn0KMDlO00T60PPKq98x+tPhV1p68jHxHvl6PWSfmRV2dWzmOsMxm2SPi2J
yM5a3Wh23Q4zLBQq1Ktxhj/BOqT8FHhyUr/t6Kjkmqtc0vjTpkdVErQMW/0dmngHAo+VNyYqSJMU
QCvMpqNa5jZzKqveKO6WEApDxi4s69qAJqqjx2qBDMSISzvlWzfSUIzA/lTmEex9aHGx7XKvt8++
NTPaKoWKV4DTpAvVHWUvAvnE9IfgHjFWpkrvGO9PFlqhx06IV4DYoZsGJqlaFeTgi3TEp+wb5YRs
y02C2lksEHXFtFjIHD2ckg+CgybokkHgmJ/Vvnq03eumoU5drNiIKcQFmP7KwKc25zPjq67CFLJq
XMZ/3bG63ltd36olIH+XfTPcAG3I3j3RpjDsj38haEcv/zaTpXecIOq1rJ5QgRr9qg46k6fhf+Vu
Rg6T0N0VG4QTGuP4cJID6MpD2Dsqv4Kx1TwJNmT8dFxCDH3H2Q61K4COAjpee/euZKN4E6zQ34yy
c3KaTK+i7z3YnoeLSBTu9cfmFDqsAlmuPAa/uIU3VlYmcW1Iwo/GSH9UMsr2hovawDY7K9aNNBYY
3mQAAuthnagdTTJlLFkqclX0kejp1ZDYbBcP3zlP9c0nvJUbH8W52BJbQd/0qmtscnheEnZEE+ee
1+dO/AZwT1gBaOPqjtqTzXqT/OSWQAvvuNokEN1q4nnQ2s944zNH+IdI6EC0OJdJgNUZ2PoY/wZL
Ri5s85bjsYTth0i0AYk6nQmMdtKVe8yrODK8ly93oqzop3zPjzD6YgRLfmDGWjI9CWZs0BppmWfH
HLcQJapY3lJ48/iJLzQs+75agJk4u/6GHESn5p0wdW+o52HFx3mRsl80xXqpPchVM4C0PhSWaTEy
c0q7dOs1tNui17W9hC0UWaAFwSEs93RU/KnmysA0vmm+N5wBZUjeR9rfiGxJIEa7OgLuO91dDLyU
nvDdg+BtUS8nJTOkt1tQvoXWIxLa2D0LLfze77EbDg+3VnR/8pLMR2M9drJbfWVcrOG8VpbAz2zC
f8uSX2khbEtEIDym4IYnU1ypAtvOfkSxD2cbXSPxi/a6LWBkdhZS3uztZKRIZJIT3Tt3C6/UfBtk
LCjwNb8Qfl3bkbGvmjUtQ0foKrQBVCeVG9PiaIJAIFmwjg+ZeJCI9F4aCYXBKjTHVDiFzhW9wbWG
GdZId47rd9Weq7l4BInmMdfRC3jQ2t0URTrnt8zJwgf0wSkuzOtwoRFKKjioeh65AihEyRX8yoIX
IUbzGjQIzCnzXRfX8uv+Rm9F0WLi+vWUA71qZADnjQiW5gpnK6q4NzIH9YTEfGPXtkS4fwxOQctP
eiRdAesosHMyonfJjv2kN9kcg/+0bqZo64cdcMSt0cz1J1k8WXStxjL6SZ6pKdzQshaL2EVIgV4r
XKEEXWaMFQ/4owicyyZujBRB4Qu0NO3GVzHaSXr9XraHswKFMUZHXX1HmgLgP43IQjyO+SJzB+IN
Rqv73wL0j5J1Bs3ibEgb/FCYyxB+FGO+v9fBiN8kC3SP8m9zfY2C0nPHzge+X2zXFNpsGnFXpc1c
hjVdy5nRsDXsptQkf/q03/g9xhGfJ0LEkW9OhcOFBJKMIlkteoslM+wotIMJaDbq7dhFNUvnY1iq
crk55G/QX9LsoDxaLyRAZpTQAEH0I+WdAAxTn/i68GJUdt8DkxaG1NBzVdWeOM/Q1OHmUqPCBlBX
dIh9tlIukLLYdcU8VguiS85GWiOoGExg81t9nwcVNk5D/tbgxD2n7SnNWQ7Fiovpv5KbLemsPB7k
a4secQOVNGS3LlX7nCt8cjDl7neRRfpFDskV8iZr5CVYSgIfcGQk6qfLNAIpZuEDOLOrxOtMUgyw
SmX1wKjd2ch7tt4+FVN5ak0PGSUkeBEgwhjZBGNvcEyjgonUPApwVV8zx8dPcDf5i4IlEkqEpu9R
ciTQ8OmglA0vzE/sSE1FJjQ45MivCz45JqcIuNRh1pq92qW/WXUicMYhr3TjtKyQtOzmfI0ppbPF
k1vBEP0bBVsyRHY/GIdakeEfGUpaTDLPHW7LuV9oYmNCcFBjrHMgJWZurHU+KQ4KbZw8U3DD22yD
nsEo5aXBWw5k8kHSjYOpwOcf8ElPk1o8J3X5mV8Ti3neheyMgMWU55Pq8c4vAktPVM3BZoQagSrg
hpKqlboUmNKcBlGTHsbZkPKabtgI2d7S5jbCghzFYCNtxSgztReCdf7T3bmIYpGsFh/zQQDR7EcK
AOGrz5I0sTbi4yNYaockIYTd1YcpAOseW4Bzt7LW70A6CbJOCIdAa4bYd4CbCN0+ZcoieySr9MgX
A9Dnt6pqkU1zjcSGMJTnPKomm2q69wk858ZXf6+P24MXPKImMs0Ch+sjMBRzqq5kuh+zJKioVCsC
kmk7qlV7PeO/yUc3DuQiEYrGs3MshUHsoqn0kwnnHsdOxwNHPHKtyWBlDeL8OxorKlMJy68ZqOCR
0h67OKTLQ5D1xtP/8iMefTSyn3xyaw8M0AkN1iIVkZvDpQnBqc5JfStDCkExTHnHBJd8SPcj+MmZ
D3II2TUE2m6YooVzJgKmIyNrfeG0dYpT7PUPs1IXxH83Mm8BdGvHslqzggSgn417TVx8rJ6JaFwR
GG8bWDJZrUthyJ80k692jeG2WfJS7zoZ2IvasGl/2aCmwd7OdtJQRDDI7A06jCufmjSl8eeLbuH6
BvJ+TQSZ5/njUMcpZD7GeENhtbEledqKIiVrQVVbIA2PHp4MShI7QGIOxKOL54MiIMHrVUVAmyA7
76hKKAJtOLeyyyXSkMMW7WWRj1A2NpOdnYC/srWINatgar+PZKgQ+R02r2CKvWCm0S1Mu+sFm1xo
huMntXpV3k70gHFgSCzFvBGYku/VfsnimQ9281WdYx76DrqCjW9Lp8yiAHdZTOVcOQvH3VdbARC/
P0KCT8emKyFa8HEEd/qVViNVupqs53v8nGIbfW3ZTN0UkdiejQsof0kW3l4p4npsc3CTqaBG0yne
ghPy2NOToMMPJdAY8j6TwL8Jqa+BwOWrBUG/Rb2V8IcQgdKinfEt7iFI3ZdfmY+ukeyQl0zYH9ZV
Qmpu+1X+G90PyCIUzsjOyaROadJiLRV4ywuLTbKhrxs1Iv/vPL5zQD2CQMy4MEMuYzAH0kudL9g5
qaXyvG9XvbYpCqgRSkNU+PTiuRMbVmmHNI260irXP4L3lF9QRiHf5bpR5kdOAyt6k6kbBobNKn7d
28kpoU+i8vGBDDikfSvI6v89ycy9Udk7a5n+odvXawD/2gpOcvDcLFCbBbOpvg06ulK6CgKGGulD
lIcPKMOMi3reiGwo6LgIRqjJssGqpQd3RbjKw9ISnEA235GbKAyQ74kS68CnzskHnbloT6dXIWd4
2dCNxX5nbnbkQePbLP6vQNOXntB57ywaoNgZj6x3fXsQpNP5XSBiGuB3KscgveDiTWlMiJtH1hE+
cQF5Vf0HOBL7LqKlZ5eS+an2u7vH60N3J/axnlSIRaJgylSVosPaXfsddVz5ySOFocrQZmvx3Lu+
hzEBB9aUwbYXv9HuRnzPEYGeEJ0TspBT5pXFnCLUwAzqfWe/jtFw/QBy+SbDvjvM8sGWeiwZTYLc
XQ7RGsf8zSk90onO4gMoIrzPftvLm5tB/2RL/Sd60u9D+M7eEevrIjkQN2djcW9apcEtHG8ss2BP
bfYe5hKT5eNiWfdvLFRyypoXj+EpktPjrwNMgDUi/giWs0ZhL8Acoe0lI+i5Chdv9pYhXAHJaGWu
HBBSTgz/iZy1D7y4SvVaF7Wy9y/pOy/aa0HA/JXWpMQps4jBi8QNpMJK0569gQjemi0uiIXjYBZg
CtE08E/UzupFLKTYTWxy1YICtDk+mgFw3SgZ/tl0xtrZSsSG2L5uAnXHvB2EqCJLI+w1OTO6L5w4
U3UEU6YKh1rTZoKk4nBe5qkDT6sD03KMb+4vi2fqTZNj8B7CbzxrLwJkfBLyT5HCYuTv0FXgbgAl
G4UIu16YrfzLszgc5/pYRVPgqC0WF6mJrEEHq9lxgXA821Vo+Zt+dQSU+O1eH8FLDe3CIqE1dWPA
4wUBU1qEaWZ1pW19rBqkSsFl1MT1Ule7ZxeFP6jPNWRdQpFgpSNrzdEbp/aOHYg7y3RZja2gci6G
aYb4rglZVQZR/xwtBBX3x3BU6M1Y6cimpE1EzMJzKRnMqw26MHU8PcZL8bO13V02prttkVU1ZrWO
NVyrc0Gj893q5U1U31aS/jXG2Ap2jmsV0zOKda+IFB6yPnNBPJu3C9HaMnX+Mb5BMRsD1MvGRUWu
fDus6tOU9o1KULCv/1va9LhqUDZlCDqia17+0tO0SOIdgNP5lIsySaJ6LAmmbHihn/KjlD91DB4l
meWjgR+qPOI/M4kMhmkSl5hRafKDI9J7Fzko87pNLKTnOKgwY+6TV+3xsRiJ4n5RwE1wlNF7+kUt
ginSfIUz0BevOCgIba5/YheMG/lwWMKNs/fBCieHlB4RCv1h7Kn6w4HXapiC/Rs53Qj7ttHixbPC
9dm6StCHyL9wNu5aZByCsEJKoFGcYLr3qTQkf0ry24EfEZZxvEPx1yT/y70h8yO0zyk7NYYwZqRX
O/6lT2RZrpt3k8Utls6bH2HdO2T79kuqq6AZvF2ajwfJim2gKOyQvTJcr8AzezsSajkpP8ivhyqx
ScnjDdtgNW9hQBS3v+oN5Adbp6apF4Ti87s6nTVxlY7dDVLm8Pml3pkF9r4L1H8+sgTS/vZWoedZ
0kL5393yqRo9/sp4qUeviYJoARrowlZAw5UIytL67tIagpjWvjSTKwFqbj3uMTbeZ/A2rSXbw68h
sdCR0v187nKdByE008Qw0y8WuaI44W/NmYe0fkmlR4Crwju8Q0oTuMSvgosTmEQcIlQyABlqPqRH
NETZnCkzDbcMa04UPcMuiz9h9byd8N1Wg1nNkd7FnzITnvCDCDooW6aV+NWoyOG+iTlmUdbCnvrF
AJfx4tDH038Kh1dmUUZ8GDzbZRa58tV3PIK9lMEIZyI4tNGzcAtggmq5410lxxToplkm8bWAX+fO
cZ3O5jx5WT7AXu+ebf+VqbdptjyWMvP+egEiT3CUX9HSeMEl1H3WUKVBSKbF2K2VhTWTr5yvBWoR
O6Od5FSzNUYsEJdC8SPGkwKYZci6OmImblfu5FXk5gNmrsUwA3u5sFwKzvvy7JwWhZkVDWe9qWmp
QyTz5ycAMNDMa7TJhlLpbGzaKRg1ImuhKktaeiTXa3fZ9YFur/HHi3VQX8f3/iSji6rLoQYtpXTG
9k9MNga0meNIMLxt2LcUfrFGCc+cxJqg1o7zGZcMAwm32oE73hibv1MB6Yz8I24uc2Smrw1WW/1D
OyvstgF+agFaC8x8roIVpBpzPpxGjKm61k32bh8H37uFNuhjnOIm48c6LEyW/GO3MvRf1UHPE2mJ
jJKQ/jSIdFhTJCmK+BRC1q+5YAA/lZ8U5T4kSiwuMmO90pJ/ifsMhh+mSsSstY8Nv1+iqaiAKdgO
qX8BDRdE537YgwCkV6bU5mywQ74lhBccyRa/82vZl4AK/gwCqLSz2uuVS1IVDgbAhdcefNXdD+Fh
iOCHo5B/+stzM5Th7Bu8ooNARM/jTRCVnObMNSBMCevHmra7fCHcFa1lbO2qgg/ByjSBEwYOc7bQ
hLKUODJSGcuQbspJwEtN4WPcHOARRi00Yggg1UqewmsVJvdAHi8otVLT9MdsX0awObesERbql1tI
LviQMZv92QaaqUv3cJlQEZL4FkdY9PK4YZGw3lBCPV4nF/xftvkrz4E9sAca9VbgaD+MsoE5aKjn
4Bx6UlhD/zd/r+dtSlTBC61KxJyO4Znng4lbKpk/7XOs34s5DqhXZoU4KdYEBR3le6HYZUIGwel8
qDuIG2EIw3LopEj9mJ+nLArWyymIJpO1IQxj9/GFlcEbhQ6YGcvCSv5hfluEfV4id0haY+fvklcs
oNDKmg3j8g5BsQL7aldgqroKqwE4M/13mEdHuJys+tYDaI2fxCKVbF8t8V4CurrMy4bMs7fqVDfR
ONQXi2tVp+NooUYPiyWbSj8P0JM6N2wgxxGrzcJCDMPWnlnYmivIqHYS49L25joYcFR9sOdD1N1q
5aP8Y9mTPiW++3fsMaUq06TOZWcv/qWE7GJyhbb58t5ixNUThzWXdgDyDjIvCv9PQ7STRwjdN4cl
nJOS6EHZqH5kidKVed6210iD8blh+4m+zZXVEoc5NthGVFVRV/fKXGlMHffJdYtKMuHpSW9duLKf
8XhFbChyaZ9Di2yAnS25ksn+/H5cm3R1hCiQcOlyjKSEKKmxJcQ/i7Ovdp40MjQlztSg+YVpoA56
Bkd9x74gxzgVAuy+tPDaM2nR3f/uPVh4gEgUc/eKM6o6qo1HDJbSEmva3IWwQIPdaogMVJrqF4RH
VM5w/S2pkCSTLuba2M+IeypetpqxnL9IKds430p3Xc/MQF3KSeuUwtCNLO+ux8XJPuyJYPpjoFQ9
BhJIBWSAOFrsCDqmX6jciBCVNV8aPlWdkJicJ+vSJin0bQaxiquM7X8wu8uuObQw6lQJGSC8lhFk
Wjoc8DktbrvXkCB3EeS0r0cSpuF4Mu5UXai0cHHlHcIYsACf6rj2w95daGa94yr1PGIH97PdgaN0
8fbokXbt8Sc4/d6gvqklgwLQAuuRBSS3cHfmnF8pKyIWg+5H7BlZwQIV8a0Yw0zRZm9pZqsmDTDr
Xp6yVrqyvWTGHzTNtAgcr7qqp7hLmVz0J7sQpiiqldVW7+Z02qp8JaBs6tHZaZ620sOcoj85lj+F
KIEg4/50ZvbL9mw6nLc4dv6qYASHNaraucU3oUBCwmZEki2lQalJDVyFuAhaDOPh2r0EV2FUxSc6
WZfY7pO12w8JmW5Ff3kCAekoi4qAaoZIx8W5pf18odQJ7ss0TbQjviXnGE1RbW902iZV+BHgW3Yx
+eVlcbmO16bOVmvoQFFwAC5cLOUNxXolJkrnN4lCGzDpO132RpshraQXPOgsPmMJQy6s24V2iZyg
8Jphw0rFRdnBaFawnrHZI5FJjXMst0GYgHAHqzklS+PX0TB3zfGTkG2SpYRZsEd8z7FT9IMZemXh
NWcBoZcyP6FuayKis9WjHzZb2wwjW3+euGcWXAoNKto2hBcdiPZfFbY8Xbzj7V9+HfYnxab84YOT
TwbVkRRTi3E3ikxTjM1gqSz8QaPkaD+QycvJEJHxBJX2NsiecKS7lCsZI/lv4CQU0ZEzxm+JGJm1
1qp34pYtky9QHa3+t+2+wK6mHaDADl8D9f7KssliPsPRsL6+b8prRMG3VpyAb//V+mpGwvK/RJcs
Rkf7j8YKmFpcgEjMauqPJq9Y34/yiXTruxAVS6a8MViSg0LCbqe1GWrRAXZ4BsF+xq148t8Yx3xh
dzn5WZU8zqLnOPoi5r5kgJpKd0N+Sd525RENLaHvO4+8EkDGDE3Q7TVfNSDWij+hUImOpiXgZvP+
INk5FOzTQRysXDh50yJA4KVodMGBp/q4Z2Qn09toP9rcru0BVnOE0WODbvZ7NasQU+tONaVWfCHM
osFiF3RtaOYu/FF1B5UAK1CvE1S2dk89ZAn2Wp6H8Pby/xDux2buMQgKW4Rmw8jAHesq0niUsL3C
WEqUXAQ7hCmXVZVcle3HbAOtH5zTrF5WcfhoZ2ojuRIt78xlyEofRSbJCIUpOVJ9gw6sbVfOnEK4
Az4cB8qVBJppM7y7UzKagMEwtxYCkBNm2sCN3r+A8nGe/AMmW2OCnis1peqq9c4dyT9cGWC7BhWd
TSBtMcIqA/leWsdIbuBY+HboPyuYIMp2ARh6LTClCcAjQfcGxbZRHhvijGbNlcqzNBKpqFKMwy57
bFM3dMkzuwsBIYPH1L+xU+KQ5j113JvJ1HZGg/xJUmg/2RiA7BzWeMiarsLWPQk/pcAHFI0v+FAz
Np/kgK4cBBVk4DWNQfGmEhT4+4yeovxyVs3OIeMOxupbAdg8cR0NieLu4JZ9Sh7BcXzBlQGrrsJY
y8IpcKWaFBZ6+yZYT/ILzopq6npugAwnyVo+q6Sqwq9389fx/Rvq7f5ptcZvXuUCDTT6mhfSi/ep
AWJtr8ncixymsk/b0D788AJRTA+3BjX5AUS7RmJrt1xVjMKj5nQXtNufR6mmuZoZvWzxWEpNNysd
JMkDg+Ufe9fvzluiF7f55+JrwrO7E+EXEu51Dl5sksuQaYmRQLneSh3/3dO4V3ufox8WlaMXVG/+
O1mEKfojFsGgsNOPmRZ2qqe+W/e9AlCoLWpjrtAAby8QLl9gMFEHWLV2FDmReoTNm062r617hl8U
9PEJ4JoncFJ322DgR2V71G8ZKO7mmHPrlVpa6H23nL1F0cVkOqCyiHPEXcUOVyTqGlYVGbhB1t/V
A8ZzMGhJqBdhFaRp5XlrcI63pd1xJqjJqCUkVMWIRLDw0tC2bH74cV/TcIyuJ7GS1bzRAE71Y0Xm
IAFGFeRJEfhwjrHOn+0i9pRTIsg+8tjchJjofcVJW0Wiwphnrzz+eAYY3wV2Mkut4Vjrj2E943KI
XWVIkHkxQYQ0mb9UvpSBTvVpnw8Yw0nOWjvAGXXfSfOKIeZhDfBOL3zGyKaX/4euTckMbj5eKTZN
JaFwHm2jh0OhdXxC+UEFBeFFkb/AiOoZcDkZZB6dPJz23s28EMp48kDboeQoDgJZvZI1efPkD8IN
GvqKqBAzB1PrMn9h63S8uMWq5x6+UJitq6W2pWOE3Kz348lBNlVnHyCNtiBmtC7D1yZy1nDC8/39
uaHDfnZPs7En5UnOcLpc5X0JXOfbLhOgqlkP8uWxxhOH0VIk1gAx0jT+TAFDQCtG1EgzKIyg2loT
qVEzNfmMamw+uiSZOJ8V1adhJwvgYJo7MWiWloPZ0C4heIOXlaVUYjaGIyozn8PVx8dE3MUD364f
rLliF1ANAW3nmuBRseGUAcKggUeAxlKmhPnACjgZd+ywcNOb+VM6IkEwdkJZeRqVOn3xHAkkFIaS
54j/MTMoD5ARj01427T5mTeQhtg8ejWDfKqlUe7dZkYAyH64jd48qRwQY+MG4vE5GldeV6vM4CDh
MrYAswlia/2rz8NZJYONSRYGq1gmCjx+xg6SicdpxD6LXE41xi7tX+BEH+luvZPCPSLA9iD89Z34
cCjG9XD6MUeA9HSgT9/zpzHrWwhg/BPBUT9G8/LXzDagH9waH5GUFFHaW2IQOx75Lcp40ihW+28i
esd0dGFu7z+L0oLbHkzSKR8Wj6P8LtJFbtDfyjhngcGDcsfnb+t7Es7ids3YmA1X5CYmecY0OF/N
hqyi5olYiBjM6ENExiKZTzteb8EffAGDMLB8mgS94UlwZi8KOs6YPbWh+9/xJfgtDzbZrzgLSULW
5T8TfpWdpJtbTam3QRMl0LPRXdKNoE1Oifn98ni4FOYhCIh1EzfzV4XrTo7jFe9wuJG2loIzRHAd
Q8B1sUZ5TQH7A86GmvHe8RrfUAV9WNO2IarqVU611CPKUAQ9sbIZlWTiIobbX4oUFC+a3cEwsaZ8
Wp6LZI/AhutEth1MBJNJYJqZMQJclJep4U+MJTmBTzCg8FB2ycBrsTvEeHqVIlKHQGMCI0mftbO9
agO5zI4G1xkBn2pqUUbYairkZfPMjj2u5fTlX6Z5z+OTRh3FQ11ZG63meXKZz+VQ2Ry4EA6TRXPr
mcx5Hj9x4GaDoWi7vaPgtZpyyJTkj6XxBWMSynDX0jek/OPStzS8UAq+M1wXOr2jy/KUKg34Xefj
cFbVJHJEggq6LqARU+MSMMg7Mq827BzWCahMqahW7rVg1WbSZGz0+dchRoUEUueU3rjE1yHg5lT9
M87dC89++EAfX6ZxjcBGc9qD4o961k+0xJaQ0PqXiyaTBLG+WEvIHMA73T35Ci9e3oRilYrW1GoG
JcZoZFDP9A7V4Qhck5C4qxavwdxx+rcG7b6/zTkrRaGfYyUoCbbi+FpCE6GNe8Hlw/Tjdrg7sPsl
DSsJyqNvoX+Zc5RW1P8FFk4+402RVKAzZ2GGCF/Zd1qeuM1rFUoTLAgze9Zn2ZkzYkMiTZvAE2ZP
D/gCNQmYG9fd9MdjQTpg2e+v5BVF9E3nDeBhhM4rsUiVYCNl+WEhbMrp+WJwK1AlQpEok6eTMxjC
bHbzBV09FXHPuzaaVhOoDzSPlqgXeaMH+XdrbIeDi+XGhxwL2RzJJt74ZUv4KR033srLCWrHyRRf
dLfuyFsKmp5ZfBKb2LImpdqMR0zjdvRgIgHU3ltQmdyrXvqvNWUZLWfbdjIanXwn6HbfWQ4h8NUr
GsynNaNncLSr+iMaPPNLvJwgGOJgcg7fOZcDZdcbe53FZcvklN0d9oLsIu2JRc2hqmF9clLjYM2i
TP73MqyP0FwRszkdcM14Re0zEbj76X62amiAOP4KGrfTchFeDEbs9rjvP2AQ38y9VZSB15FZBbKO
O366HD5Th2ITO9keyK4FE/i4/5ref7kviMAU8yasGAliC4GT4OADmzNohbPGYjUzmXFbVSBJC3xv
exLt+/uw9FOuYHj3TLir8EhtsV2lyUkKcb+8TZRxUV1CTOs/s+KaddMbLTLY6w+E7UIV8Ko7iLpP
J0mvFc38bhOFscXMekHyKtIxLM6wuhrwV1X+ZukIYizmO9w/VHHztqkeBzq1IwDv5RAkfGN81a1V
OvfnOFLdLkjCpAt3aEonIRTDcSA/iC21XQPjnGmud9AB9qxf3m7eXuhgiEyWqV0+xwgwKSpgwU1b
Ha0zHTFihUmWt7WT4VAU8W3ZJM4bIuALWXA3yt0zpj8CKFq6X7AfHUDsFliQPnULtK2mVo9EostG
kYpOuV7/Vox/rJrMBKIUmCeEIe2D8b77/oIWcrADyCbMFqOCZ6mX3y8MjojlYZGvBp75rWUlCkO6
8Gyx6tSKfDCnow1lXMfAueYCjPQUWGud8oECbWV2BE2yFRL0TeieAM5kgwNBHP0Wlcr15mvc9IPe
ULZTR7b4pjxkHi0rSm6zYgT3thGTFgNQrBClFOhSpgM8wZins5iWLY91EMS1CJSPl+M5/PJls2Yr
gyzMe6BQHp3Z1S5mi7Gfo0ZXS6ahN/KKe3412fdOsIXCrFoU/KRFxU6ECk4M+gS/9ecZmc+akzA4
AB6Hskw/DZLcwRrBHOnxiOEOJL7un6F94t7sV1bUcYimTQlyaYROWFWhZNxTkz4A98EKVpo2j6+h
Jvz2iXrCw8WqbocIwJj/UUA+xIKzjM5dfOyGIHDbDyhb5TzgZJ5PqsldY0pqeBtjIsyE17UESQkL
wgH2vo2rs25jVs+srBbU0vCkg+4PF8rdIbkRW8jAd7b6r5JyrziOXw3Y0rKmMRHEpSkZ5WQHyU86
GQH0VzSxDd+0P4qJaDND1g0g/77LlS+OtsxJT7N4IhNUf/6EbfqfTq8vI83PI1B/yG5XhlZlnFRU
KrZ65KuieZiS5k6CDaFfz5FD8Si02V7/8jPuqcM/cNEy7DeMJah6guv2jq1m8XYRbKe5hpUD+cuN
JSVRNEBM8kO4VpU8E4D504Oa3KNNa0jI9a7Wfieg/B/U11MKrExV3nu43vApGqYlHcxMZoBVG0OZ
6iAa92t0LaeeShbXpbzoLKPiYBwaOhQmj0qj5+8+7o9fw3csq7DLSjmIHO1zoSEBb2ndJc6KAW74
8gpEwfjWqZKPKeS08qVgR3hqQdYXHKaTx2S3OTM2MIEnWu1TzNzFOgexkKItI0OqxKSx1prZko32
tA0Qr5dya2V+XsSQDb9lg0Iag7EaAhPAhykuv23xcbu12AFlml+LczrN+XIhzsBiGnxUmQlIa/8K
FwMVpRAe6AHjCRx2WzSBAR/i6gCpt6/hBaLjZZYzXfCuE3pdfsXBw9o/GIu+4eYEIeRzvsxcPF39
Y+fQ2do8vg/7bTTN27LNFkWm2HKjbCDQSOa8wvYNvyJj9EIkkuAneavUei4RrxnCLzi+m/vhKZbc
kh+lxX1rsbMfkBWjlAv/YqAko0WB1kkFZJIG2oJAzfYsHagmlauA4I/lRynF4OxpQsu8+KRhOF6U
dhxw7eH7v+Vmi0bSmishXrewOoHt7JWhXQ/wx8RMzXbd5OW8u18eGgNi34DODLLBDuX/71QUhUyq
2zuwHSxa9+jdPRVaxq20RaExCkyz/tyJut7vWvYhMpDW8JBtgUtFMAPMteOskfnVRmNh/9Vg8A+K
APVq5phcId7yuB9wJ4vNGrl0oYXCns6MuuFAtxInyUAn+CylFQJ49eJ5hu3Bg8mSHmo9M4i0IlHn
1Uc9Rr/OMe8AB4ieriWi81z1g7GsPGVDvP6fna4CwOvvTnFKeIu9z1iJ8StPcAK0lfIePd+WF8Ab
Y4hsi0aIaSa8VzVSswwE6I1z8RR/Kg5BgbdxKwOWkSCPqi6+Ux/L24rkEnZcucWwuYpQVc/8zUBt
5CAD6tPhlkNpXlrs4pDMAKq239+V5SPiWYGzeg61DtaWBb6KLdcCVp36XF+lXraRdBqq9kbgQ72K
45zwAZZk/E2PPjk8796bNFPDGVp3TU/ihQQHD4pHicDQ3+J4YdBxHNWxCQDuyCN7MDqYTJgBZdLA
9K/bFc0VvaXLIvt0PXGVc8pAoSnmQ6Fo77Z6sv3Eg1gYRRk8wbEDuAMGumMxc3Mr5Mwq1ClQ146C
sEKmcXE4pA57wH6rWe9xp8x2AUDDZ1G+kTDa4w7h4CVQv7cgVtznKTg5y51089I6HJmpWUMmWlAn
94Mw46jJHP1+sm6L0sSVs+p7yvu5BS4MX7uXXvJY9LXsXfYJKqGni7C9PQCiNwiG0tRg2MECGHPS
WoUtyOf4SpJfc6pJnq+GdNdS077DcJM9OEQ6RPt2pi/QSlWQw9CW2qSilw101hKia3IVb+6yk3OP
aLY/fCpVmCUEmDZzAckhrGD+qH5Z247J6Fr8r8OJiHPwbFuYJS2eTQwYsMJbBHwtfd/LOpfO8GNa
Za6/2RWCP4uwQ1+EgPBLIQGiqD+TCWV+H2EnO6ebVkQ97zi/NntlIMm6OxQwrBmhGWNmF0lgwdap
UMZlJ3LF9dnxXFEwwO8b1/JuYNd10s0mRMgqp/RS+pl+Jc2flnkfBfEqNe0rVMtfgXoBkrQZGf+q
yfubYMDIDEHfBE4gROyhj5pMqy6+LWazizl49oL3Qh99u7ZpMiRA5UsA3+7DRXuAvjP/Va+4jbhz
KzSzbzdC98Ifv0TJkKxjC9QSAqcMxx0ONQZK4UYwOOVcQlttKuP7lcAkHHbdPsUgY/UTjwH+ksdE
L1A8g9wVvEKzNH98Uc+toGgalkepvQ917LYkx7WkMXHseNTcDr/ned9tUIr33jVWJORCQAd2yZEb
Sk/ISku9vY/dlxNQ1HXd/atFivbvcyYdKUOPw18+L/IE7RmrNyohplBWTpLdjxzGHKlpWwmEStZy
gRCXh0R+okSC6DOa3LexYo2VNSS02tXQqmwrw6jXkxsSaOsnnc3DR8cNGulTB3IBoXfk5uk3ovQ7
OkLVtUL3pp8RCfs27QzxYMbhMsgUC47AU5O8aJEbYB/FG51v+Lqj6KJuD4mIK1RwMUVFkosmXFFy
krb58nNpZ43mLnGBwPnfjpLEjvkUojJXF0fHrer28m0+vVa7plvG0PtGySpiL6zzkddCaAizdNpT
x86vJAXE1L7xgS6KKyAu6Is8U68grY1eDfmRh1mnh7DIio32C5U1DlPJ27131fRtBatFlQ4E9vRf
7CyIYjJdFYcqddTVJmOBAYIqBtHJXtBfX2kw+UKGP40h/Ry7pnTNlreTNb9aIIZgevIplMT0ZQPf
6YrAmGeK9byy2a6ELheLUwKXFXYuKqgL/D2BD2KHFy5jbDR2cO2e64YgT7sxYs4ORzRkQ8ybfIVJ
KNyvjputI+2XOYSeVO1Du07PoasHBGwlRSoO2yZCbjdPlfwoTmlK8wXHKZm/C9tUoFre+jThYYeN
JWLIdgqN4oLm0Nfj7KAlLgb8HbPiTP96ON5oln4BAwfLTmxzP0bbqLFBWJYRHunJg4Engg27Pcy3
7Ky21I0N/BabRxHPsKrGoLxb3MWYudbhCG1YDu2JyKuSkeR7qqEL610vmg9m+JbV9skn98gx4Zpi
glIocZjVL9XLv7L8UF8/eHf2yphQsMg4dvlksXY+/li2qRWdU3avgC61KXknE9Fs31C1LwTrn0y6
1Oe8qbFedMwH1dLMsJdYWqfBbLXd8gc9GuX4iyjnsgCvwbhgVWzjIaWMIZFzVQbyVKp9+2Y+DcEH
F80c/bV1XGRCE9UNocm21lRmB8HzHr6mYeelxmKffpkC4BP+r1RuozICGF6nPPb5R6oHVNfmayVC
KEDapuI1LNX0sJA7emm1JhOW0UkEUDwGsf46Dak/Epz6uGsWy1FNzGkgFbBGCFZ1UnseJ61kPOaM
j/RRXTtwNV3tbzT29e9Dz6GenuUeDX9/CNf460Qe+IpRW6hh2sO3Mbhr5qfja8/lIZ8RUdGXF8l8
qG9Jf44XXsYpPVG/hj6cCUkKntvwxZd1WEwlwp3ZyTsSAs1LK+kBcTYGlQGi/9CpCcJ5jucCYqt1
7eUGfwheUVXDq4pf6Lvct2IH2vBG6cQ9/Bke7TEu2lFLIz2c7sI8r0e1rdu86OAtMlpEMoONUjP1
RVAWMkC94sRRY+NorgSJKrrmSzKlhhuKV9uSQOH3ui/eqNt88CoJw/+WUZE5L6zOWfL84KKJ658J
M1sutBHC2LoLHDlqowmRiWqHyTabFLnhZ2dpQ4vevdB4qW7wK9L1zOERsn+qVc9DgqJKP6Ob1Vbg
eGEL6+URjhgVxXO1yT0C4NOdWOLd3EZn1ugUsACMXd86E4u0dLPTNIt3iYxarFarhdL+zWJahWyH
DSfnFuro+urGXE4C9MjibIA7qWoEiX1h16tYQ8FIYP3sPImaFtTiVcrhxP5zPxIGPL4EE/yP/Ayg
aVogE+DOrHgrL02AxTG3ToUhzDdEegw6NI6nWjZmKKAtnY1jP1ZAEZUzAsSkiBhqGCCgGUxjeU99
xNq1NYgq8bQ5z9il7STy6ULpDcG/ch9HJXs6IzjgAKbdtRuDVbBH53uloJP6BIf8u+BgXih29KNg
70TLNPEq6efX6co5rwUN9oeoEPaLJEeYIS4uHw9lKpuzHREpraw0Bf2p9whkrffMmb4KN8dQGZnD
Z2sVHPm/o+Fe534iRhCtiFIlbxYanP4UYqiuk0dWz7rhutqWVT4oPb66KibkAzyv2oJoHvRA7Go7
8K6b43nx/h2RundGVgSaNWwtm6CdaaZjW4ob1zkC0mIOhVq++NQzS3kSZ8PaqTZVTaLy+3R486vH
So8rVb3UXgn5a6jGg2nWK+7a0LPsPhaVMoCplmldsMY8VH60e4RL4m7QeU3teJ5gvhiBNH1OZhql
xPluLj8x8x4HKN8YYpYeWTrot9YZT/X5A0auAsv9SqqaE1yuDo4xujXNueMBJTfS2EbtBUPWhIEW
/PLiV9Z9gc1onkE72Pbg0cPBKbZXI7NUPDrmbgex3gN6HFoq01yhU4Mwx75kOs1MEHlgDsD5nyyY
L1Zug01Ngbow0Rnw2RBDdl5paBqE0BeLpmutr1rDZD0+eZ1jXHBJ80KK35PkTAycYvvZMAmQe7Un
D7aNK9OuSwK6Oi7z3dy2VaBLlGGRqpI/xxAvJcy/293lDnZIUL1cAwRbF74WYWNXHYIhCVtJJEDx
A4O7ytTxfUDrdPBjVmNoV3VBLXW0hHPXQg+LMCbtDBc6UHpY8xL+acndpbvdpaCBK9w7WKxKtkNW
cM/ofK1HuOUnG+QR7JyAHrOuWV2q79aiwOiItoZLRrceFIUKP5Q1cgHy1wSiKmkYJjGI/E8d1xS8
oNvDsyc3U/q0zn/gutE6zBaV2+uI6kQP3LpI078c294B4xi/We3K+J8b98HcAgrD1aF1gJAYA5Ax
snLpFWxu2IMZriU8g15YTJHDmnZKB1IBk+vbloPNS56OCBX/SICTPzzf5mDx94ry5LlPIheWcQXk
tYM/xNaKzgLalmjV9MuXwm5OHInjNBOM4SYXkVcbwHiQywDR8ujp+vmozBD522ObLlnQDtyEw2yK
zmI4JrWNl3A40jWKYl369f/VzODS+AysvST8R+Hi6q+spPoYxJqt+sREEV9EZ4awKQzTw6tae0V1
XxQ3Orgu1Gf5cNQjNskVIEgXgDQgM9d3cq49j5DAw/Wv+Ho52i2vFlq3i7Zaghq62yv7Q7FtD7oR
vg3bxxXYUd/pWmgbcel22l67On3bC8Zg21/DK/R1aEAI5Hr3nFoWufIOjt8irPX/sKLNQZplhpzQ
wtfP6for+pGR4e4wOUBIyR7BIfgThtd7nt+9I06GMZcfJv4s8kGNhIZQWokugKJAIVGc/QNnFU63
BwHW4LFRevtmgEapAmiKc9EHgmFLpQ2N6CMxjrmGewXsIWl9JQFtb6bDzliN3R3STH1vI5l29BeY
CSHMWGyjGcLxJwkm/smcv2MhC+kSyFmuf8BEsA3PBMxJsF6JA+m6Qj4GWVwCWUGqkO3MRHzeD6QB
EhOpG/fCwpykRarhQlSOGs4tMOIgokfldDwLFpAYwMto4ctgqdVZ8PGfOS+0VbAMvulIHRMfvx2U
PkdvpfNfPJCnsjituAMlLhQ8TXFTweMBZ58rnvkrAY0LPQa+Pi3a1a8jSu1UEnpAy+ydIV00WneN
NB4CnTLqnPqfpNpcOZD+5B7R/fgS50QqSW/Fjw9+Grpk52RlFDMAIJ5LY4IaSOSnQCAJeJz2wbRT
A3YfdO+NkB2KV0anWgo1bKbjGXjhZYq1pE5xhzci7DbPbm6l0NKQQIiAWS1Fv5CmVx5BbhBROY3V
ZeLDF9iZOkkviR+EhaNJvp2TB+VVCTqAHKB7jsxKY2COXw2mm+l5BFX7XLN5dUpLl4agjIjZVMj1
gBczotWqbUfgNTpp7qM6NBFc1apeZbWTFTYss9sPf1kgsDkVz/ex+ocjWAXG1Zr3it3Ac2MPAUF0
OteqMOmCAUkn8deqyYbrM8iFQjLyuKmdLOdhFDsqOteA980/NopQkQZM14xG720Ly73+TLb+uPR0
a4jokZ5a+XCBaISikPTkTMFj9EtRzpuy29h8iMWBHZAX/oHWmqNCZ3OZNyHXZWL0rnTIBtDngFDe
tmp1JhKbUke8II6wmluU+uRSalQb4kBHMCIDp0Rg5yQmNl2roJxO5pE5FiwpVbci7JPUXGzFij4N
k7oBp2ZWFRBy86wWxZMNEk9wTTiHZVdqhKHn1zECWDyDDa/qWoPdFbP1A+ZRaKn1l5LhJFWrhejH
z6omObUS6lPsSyFoauUgfZc23RuOwtLmB+r+DrO/rQrKwEmV2x0gjBk55uHFYECjP2n8fHusl1j9
2PSyVwDM00JG/LMORhRM7doZjCGYCuoibNOy58z3WioWwlMKcGiizmh0AKRDgiKJmrCgcO97OVq4
0N9He8y0RoT4FXxf+lSzpSDMA44maKvGRkj4L0UAT/5j8kD3S5QfxONQPl4em58rZXYZg/dHiwmP
Qjp66+o9Y36+0/gsPt85iA1ewrl6dTalKU7K19jw1ofucaKXjQBwoW8HhkD+SyLy2WTyD6brZFBK
k4JaM336uCD5G9pkIpUXP3BuJkrHv8uNX7rEZ6Q059fygnuDgZfbKeYr4buXyUNmtFETQVpx00Yk
4x5HIPdb9v6yL531KkOHfdtbP+LqIDwBvw3ailjswyQXMGhHX1ZSSijskS26asDwTVDsCXkB4bYs
NAScXu3+O8686Y/IDhUNiB9N5Ol3utPRDrd2m76t/gMijQFk5jKvDr5r7ZWIMB1axDBhc3I3xNCQ
UDXgVWImVuFJaW/wEBTuvSAClDJvnBhm3M+Tzl5opE8IsE9xIUSqXL5pPxtY29IMUTyR1xZDPJFu
HzT26vniNtg5IEv18xpT2XYeb2/mPNyZYAYqL35K9KxSdp/xn3RTCYb1PXZgTYqLaQ1BMJObX8/T
T2j+svS7e7sPEOqNHSHtzDqrP1F395qGQ9FVXW8Ha1zUOdiJPut/GEuQKqrpeJMfbVTdd/4pveuT
txd3SEJPdM75b3J47xr669cphQa3Y4kLCWx34Bc6rVMvRnaPH6IYMgxaD40SLRAjH16j8ADGoUht
jU3yuUlHzmGLbaIVtVX/PSCgk1oEVw+glDjR3GdZZIgttOvsedolydMCjBm0Harb9PtNC9pY9OvU
OpUGlxsSlzXGr0aCNg9VH6Z6XaL7XS2+tLIJpm6L6ijwzVgHzc4aryd6T41tRWDxks5RYjZBUpoC
yTd2LnVZMYGHXEkcBgqin8q8Pzcv0YMwxVsBHoHMQxdn0NbTpsef47hewWIEf+NwsdWXSo4UtWiQ
ynkH3ZLo8Jgy38CPthgrmbPVMQRsqufuL9ifC+agmulpJ4dryhfPpE/d/bietaY7Tq/nxC+LSzEM
slz6mnCqvVevSPP+HZDoPC7Tcaq6cuwTRB7skjDFbY8GKjlJRJUtITjPm2OtsWcrDlpg1Cuy6bBK
afJBJxoTXDjkwddKo03To6n3tbEHu/M31HtO7tJAXClb0BdGe41OMtEufh2gG8HFZbsRA/Gi8gGz
TIX1u9CuoPPWLAKsWXDl/8y6iVDYsY89uzQHevtO1ZXbTYV4d7JU2ZrX1t/7fqbQPebdLMdle8m4
YY1qANslVYfbnVg6E3KRo0vZ5Ctz9Jbz5o+eE4WuhTp0gVE50lNOjaOM1NzaMPBPbXxAmSSfPVlH
RIn9fEcAMtAGK58HcLLV3UIuSWPfAON6GounEX/SJAIK1fdoWmJ+COSXMmLPvYdEQ4bnhhuL0des
+XddGLzLwAffPeroINT4CRuXvCKW76A7ggYn2vxW1rWouik5CVDEpSjGcMKV+FhDh8+pUa/HHqtU
PvjEFLwAdzFN3dWHQNerXDLYqaeEvmDw6Xk3NLe1ItRB7ICWh/R7vAHCmzDUIw1tY3vtGrPF7RmY
9zptriGwXbjmyxt29PUVtqypZDipoHyId1NpZRnjSIMN2K8aHvUotWGUrZwK+6TIN+2ocuo/VoS3
cFl49H/XpUKnH25vtDNhrW/F1mo7H/ov2f003Hw+c5WTI46P4H9QzIytL2BC95Y6Txzqzl6DnEhw
ZQC4dRU/RejzEQZ8f31PwldkKgKJI7mN0DqGHTcwPO1YXSyxzI2nkKP8OGISAcuuJz8ME6r5XB8s
5WwY67zqijYO4fKg2CCpIj9LaML/Lq3Or/0KJFItXieL7/RWu/+Ff1C2k+DTIRXH7m+uFp9Wr/+u
CjIG1+LRKxv4L5+sZJoinm7bj8bPS7GSY1FiT9oNuo/jgdBLNoVbZ18WRJD8740WpUubOk2KZfbO
+GGXp7W8eZGpRiYX0Eo2k1fzjDr6KOfoIBiNTyMs70o+ogf4AbkW1PY76XPNbie0pe43RUphA1iN
ANKecX5l9i+/gMVJFA9w/YOOxYeeuVM8EUhEDKoXXqTCEJ8RGTMn4VxxNqmB4d2Nsn7uwRablDH9
5W6iV1i/2iKXu/tA3K43R7mn+8HZRtD+ebGtOqOStvagSmjfRb0ATddYzS3oGflz46Uv5b77gvGh
YEQtFqRpZ28z9k91+1gW9LXSbc1NrAoDzALyFYaPWL1qvY4aR9l/zY3tW35WmO3mjQIJxaR8oftM
9QoCuPAhEwQFxvzvGu1kCY4Qazv1aINjy5jCeO5a8zbNBTlG7mV9ualonsNalkkbTVYy8Qw/3ly9
fZ0+75N/rk/yqq+bDeyKcqtr+Xah3B6wRSN97iGgrgG5xQ6XLH2Saq7sQuszu0PFscoW36E3THbO
IVFmAhZUjjWA5oib7NUosGrlpE6pp1RJ2TFZ44gAdwLkyNEHOSiYe4vT1HxA1T+AmJQCw7hL56nM
G1kHkvVRdQzONAKfmKUWEaFF8JMdc5YPhhuXeyik32SeKYLZ+U2PP72YvEACy9U2k30cKqWKzd2N
Nz/wvIOOQlQYQXGg1y15GZUd8mNu4qVK5V+qC1LNYgwHGc0/+K3P34dBazo9R6WFpQyfhav5AHNx
3xupNnT3VwuEqUc2DQJ98uEGrC2h/KCN/cz+nuSUvPvHgocVmRSH5jg8DtnTgv2Z12ku4h/xtPRE
CQtpI0bQxwLeMCJoclv9ajX0SimaL8eH7wYI+n8KO6vq6sZ4EWztBXidzPV5EP5iNjajIucgodnh
VPo+FxY127VU1NqXGXXfjVqXJNbPO8Q2/yAYDjeLKiqivm7nPa7eDfAD7gDDXdW4aLCxGvY7fIsf
euFYbW0QsujCoy1n9KVWPtWfWPezXQWYyeFSJ1zmir1tisQnFM28s8MWyXP3dkh1aQN7hLGuPTQJ
jwSa1HTwcpRpFLWacz6F5oquTc8GJcAcGpVzzr+lV0EZXqKtSMCswAGSR1Mf8ZTvgN1nqSsVp21G
rA1ozRsdf7cvI75AHSlkckrUT0OhChoxrZaoE7VVxdIMMBH2W/HNV+U9U7pYQTynvNF3mYaGXCs1
ey1vAju6kq6Tgbx24YruqKxkR7vv9g7pFwfy02IspFUV8tTLgAWu9u+nmoQKMlMhb8wAw9YNLB0p
ZB0edS9W/W8TkEkIa6qHNoY1dCay40TfC9mwA6ETquSHN1RJRJzdR1dT4EesHmxPkqnmikDuoLn8
1xYTcNjXGPhJGIyBIWUeSAnBJvTjfJyUAYRKPC/CFYo3j58GPIIJTOKt88EMVedJvJJj5pHWJm2+
UXyGx9tEQR0cV7FPrmm6LsV/UHhsMiPJFS5zrHs2zuThDO2Lbt65pEJiqRBWUYG1Tnv1bQoNRu2O
h1XxGWwhXKu/wPCWsree0Pb2TWnyX3g1f2vY7pA9cSK1No6XlLNl0nx2SOiJJQ9ppMyFYvjmR7OJ
55KBRbsqEjPBI+GAdX4UtH9ZXGFABM2YP+TPL/8/ufHg+lX0NeabZB1zfLoj8SEdGcTuNjOsP/oz
xmLTA8UEcv/da1KiQGEAG5MeuwFoZc8DFT4h630EgwH2EB6KuRQOG33IPK9ywi1NWzvDVcXMR9d9
YFaEoQjQwVklIH0xy85zC0QONnOkxjmQHkRibsykVMa1AQy5cG+4498m+NCQBHBker+Rvd76Vvi8
XSgjEvyk0HuWnhjX+cyVeRjsXsZM7c0ozOQNSERQ8he2isAPc/L03WrkdxqdjGRGvYpp0IAtwopW
f1xhB5d9OL583Z7KxA63LCIdM+RRZNpn8dqL59uZUIuiVHC/eIUyMO6OJ9bh7dYYJ9umB3txp2/B
/w1kSBuJnc4rgBeTGcW9A3lmiitesE1UnzO1Nv6HIVOxgROZXKuI4JJK9e8C7c19Ds8+9tVcErtP
YJWdB3SYku9avPbwDP8hAF2jsROZzH3dXgwC2v8UPrm0F0F0c9iMKYG2QeeLh6/jmITAcjDGMrY6
tRLoOEgRhr2Xbtv5tAkwUpK7dmXRn9ESszhssjh9qstk7ROMQbrZhG/ypjLjrHIa98KmQKz1huoE
ay6yLuvDtVQqWLXhLECVVOuzwR4VtWr5JVTIDD2B6fli8Db9mMVdMWEd7sozswQwD5wVppA+mIXr
aXSyJzhSQq0lYpHDAWegLNUADDXaX9HBnqL+J2pAVyLYhcSD9yv8WHWTShXc0R4Mo0uok04ALX0x
M0FHzAXGBD2eIg8iyc6EFYxzv2+j5e5Z7RbB3SBlJHpSs3qWaabmbN/XT0wfMAKpfHz81HmD6Usc
2VGZbfj0T4T0yP5QAceB5VqJoqmHDJP2ClZHU+FA+lKMXvLyC4xEOjvpWiYE2NFiHMJXg2sXWTUc
jn1hvV+x867/2Y/hnF+YcmHSzrbiENn2VCgPhp8UPJ7XEmMVNT9B/zKsXD500FdvRsTnNIo0rtgl
z60NEffgcVp283M1h9LpX9sog4dRjAmiPwgsEr/cTPNGSA8wpuB7MF1g6T/ykr1r35dAMqjf8nNF
9QqeytUsdxYpksH9UqoT9MiNAESr3gQPTOd+cippxxXaL07nlw3uzEQhmINTabESE4Imo1xjDLdC
4CJ9eD4Q793SIUHYTiDfofPAd4FY1r+97Uyagm48r/ZQGAftfcCUgcFx8ZlRrCPpd2sqQge5zyJG
dwqq3++bSJ7N9o23pHiWNZNj5KwVNsxj+xDg6KK0mG0lpTI16rbD/TE9K70LiehhfcSkUdU4jmU1
xit4nH+Ma+9fJZlJV6MekMn5OlEa5VkzRfEQK3vJXrwOgkpWXfkG/Al8fwQQKe2cRjwKSORHqCUg
H6KPR6pjllFBcG1tjK4HfvZ/+lzRfvtqPtlkW39AuRtikO3L3BM9y3pol5Tkx4J1G7QZW178hiNX
4/lXwzgENstdqkrgP2qCwnNXFpjn1HUQa66uVCpev+i5qlod90x8AbRGdRabRlIfBSr+0Haxohcu
9wwU2h30ot8ibhsi0dsGwD/QZ8jf+jKHvVjZ9N45Dha4DRACJoqfH3UccRN+WZoOe+XkDYO+bYXH
OanTVZ81d86Gnxv8XwOPbiSIQWJXuz27HbbAvFsrMAWWXiW4kr5M5kWZI46+0C8idE4k9O23N2A5
CVsnqd9hZneNGAaXei96+BmgHvCIRfpMdJNNqi6WHbSo7ZVGF8WqMl7Jq47cJRG920qDD2rZqQMt
2y0LDNJZua1IxXx8EeLWmGu9DfgCdSClO43NfZA6YnN4hM4bw0rmy/wg0YANKAV+wO7ZrdIiErEH
Mgn5F8uL2+JfFB+P6jzEc+pa39Xu7m/EsWClQXMDK8+P/SDcz5f8Aej0CiiRA2kzcU/uOCNqI2Wg
zvyDx+cKO9N4D+MHstxxCkCVS9cKVy8wttU65ItoBD02e2+BgzrC8DVG1YF/sCp0WPOBrKgOVj/9
LhUGaT+aIQrEOuh/ScLg4GB/ohJDm/58csXPrf6/QtJ/2AkvfwC8szK6Sp2p7CnHRFizWoUwdRRs
JPvysasbSshsLUsfUpl4tmlPUkOAmyFwkVgkeJcL62xq1+6rQzFXWYo7iawyY2oHJYawe/+hpbNa
qYBP4ouprln47RUf/p5cDfiO6JDEIWVybtiPGhXTAvygNiQTapIzedkLUB5pwlPvTze9RVNo4ckQ
aoqmLft86zzuBuhPRgX6wBGblcYMJ+d5gFJe7TxVb2a29O5O0FvW0i/lRGX1JlK6p5Nfsd1szkBU
9bbWC88pryqyV/uUR8WRy2bVv0YggeGuTNoowZ99dU2auN4xps2QccpM2TnZA0KFAPXL1O8QbxQe
H1jNlqL5J45F7to0gvr5Ka8Wb941YtPbPulPmCdpX3eYswtsMbbgCPNamy+tCw8K0dWEKEEWI5Ct
4X7V0KrasF6XbMAn424q4NB5tpGHvG/9MqTl92Do1YyfmSe9itrD6zykvN+v4ZYDGTOXO69ROuww
NDYYBPMeE2huXqb944BUe8uafuHeXbmlx/vgh3P3zLrVcA3o393Kv178ZLUCOwWbCsAcSaPBNeH2
KmhvWeHsA8SeZp0xGgXCZd9aYxZL2R1k0kpcXzOLtE61vAa0I+p+jHwOv9jTW3F5TxokOfWiWwHo
GHOSlGy4brgPzJDVe8C0Mn/yvrh/n8ATYRIbRYsSjd23a/JiCZckWVk3Et01x7WRJICgPfGaTSTY
QV0q9rHaQnwCLeJoSRNnFTX/D3NN2oxfTn2Xa+gcHGiL5YOL8xCHJeZEXHqvis+KJOoviiK4UyAI
6bUUUIl9Pt6E2P6SegXAM/ggKLdW3oZSjVJNNwAxCRybbHtoIbYH7JQHAROMKxF9bcwkY7szvsn5
uOJI20LThzDjbiv1qG7zr3HT3iibNwClSP2Um2iGHWhmBYHcyQcN7bl3ihzxa/Q55MK17k9Hj/mf
LDUC1yOx6WtuL01AI7AZdvCx79+66K38rbuxY89auklOlYqndPWTjho+FDTY4yDt9Rdgyyd4qIAR
hVrUt91DnPtmob/dsT/F8JZ5h5du/ZirEs77SeGjA39ktvh4E6PHmMp3w9sVOKnet/281wnmBrVi
IP6yaWLswO8rYM6RH2ZsY7YXbJD5jgC9q3kSZ4bA3YHTer4y5zJyJxM1vc5gdHkPRpWTF8w/CLtp
ugU02QjkjbtgyvnYo70DA2lEf24e985toQd9qj+GENKpzIRh+Mwy21Xqazu6T/2In5MfzjYdqRrk
ZHhXM6yDqNAaGpBnov/VgJorH/t0WFLdLtFwd1rWmoXGFYC2/f3U4uhcmOj9M4qKXqmaDotJVtaS
0eu81Ry2HKGNT+VeIJ+6XP4LXljGlGu30Uy/TPy8TPWka9tp8AkmNJP5HCZvBgSW0K8mR6FXv+OQ
V8k3mbHIA7OZ6ooFuwE2Ji9nHGKS8V5nFEZTVEvy3GT3OONaepry4ibvhnrXC8di1HIiL4Yy+z9g
kB9sztg56XQy6M5yQW1EAsYmFjyjeQlVgxMpYSqJKuecHgKnMYEhjkljWXsmFRrmTEZVFAI1vpRM
1l/Wb02eo2NO/v/uX7gW5GbciOVPgPE159sUpMJQUqIaNueOYxq/HTxpyFn8I63Zo/vJ5+HZBoYE
Xq2PCSQFSDvhXkEQQI8RD4Lu681Y+xKEU+erp+Sf+DNUniRq5KpE9NgegJsrwkFEawbRZb4oOsY4
r80tYxgG+lCzz/T9gpTmtcknL0f2xPIZbgRwqQ2/MGf0bf6VYY79+o3AzIzlt9mmn7oNQ6qpLQF4
GuTDr7S87CKUFgc4B9bzBVzVVHzz8VqSxmfrLJQy/eojd5eKPfvMx37gkcUsEFJU57E4n0DcWCn5
+mP8R7YaH+BgrfZkG/5XAaRBi6cRWgeegWc40pIswyN0+Q8kWqv3MzvmEFxm//8XzLsFYw0pThNo
MHDqkqLUQGcOblS8gQBgDQhMFaYX6CEL/iHQyWWV5SCE1uZa8svQXr8KlzXMYnR14fGETBLrbLl4
I6I2yRo3JoV/qhPKIUo/q+HQ2Rw0FwSxNLiuzW7moGqd7o+QDCQ/na1WcC6y+02xgZQq48NrOlru
Wpa4k4Xx6+bI74nQ8ScbJHKedXvqNtGD6HW3fZ1LDMl43gpK1I58IMcKSvCj89TbVJFXQ+I4YmCA
y+OwXy3WGrYmxWH4v0BAYvhPUTJKeIN1Ow4Xh/EXLrklh62Od70VqtC4fXxC9Yx2/vqgNoHeoVbq
QmkdVdA8yLBsvZ1kwMdEA/R29hxLkdOzRVdcFtk5Bh0MDzWlljXp4uQiqpI34Cx2NEB0uTkl2T6l
cB5OxSdJK6vIivrrdXsxg4luEjVCp/Ka1+tdbAUfYm/6/w0aeEBQ8owQaf0rJr6i77kZ3HY3PIg/
LDhSq/3NM9PRZAi3oWgXpcz0eaInq0o56A1w0/es5CwpRSEhknFX5/7HqXso3kIhcixPE1EDOj/3
5S6LNNJVoPW5jFJFqkhjEe1efDaB1qOnEgIsT4RXGrZyeMlDoeajsOwnpVZQ3jaOQ3Iwzf7vVb1s
bRvCs4onQb1UFx9kWV/twU6BCnaxK00F5p4Ns0G11iaIb8dzUQ3yx1F1fiH7H9nm6kq0t3rfxt0D
jWZArv4oVNyfk6rEm3ExdSv2VgY19rWOodMUOiP8xctGglFg1g0sj+FWpU6Lnab6eUAKoAAFfTbh
ro9QByMItxkS40TfyhWZrUBOAKgmpKYjAAbVBOZiE6uFGkrxZU7swGE+Yu4pLmhvL0hufaSqZHW9
qjoiQOx3ihGOE3CqOKUkc13j91wHWahmkk2lQbzhwBwsPfbsOdrmkLOMla565QLZzK2xyXNp9T5y
fdU7eOKe9894uRl7BVwL5c21MtYzHdPoApSlGBfF0NIK5fPpUVMZz0vWBd+INYTcfH7A1UY01g1S
rIlNbwf2KvBnH+kXruPqxbKRIuPmPx7eICtRFVXuWOzohbS4wSxOzgJolALoi/0hyjth8JpGQmd1
RCpdXujKfqquzdQSjq86MrjJ9LimyQRNgayKGcNSjPPUZ3VSLYgrBt/nrYtQcn5L5CS4iaMoY2TI
odsKQ0iknLtBDGzmmd63dwrXX6mZIq+mDktZcYH0N8X96bCdIm9w3PSn8Exjpk365jaB564i54if
c9op89wWj0ePIpMMnZ/0no3ZstmOA18hfXr7mMzfctYreZaqJMJKvCq5UpU6dOpGlul6j5j9qg3G
I6OqLTtBEPea4oBsaaKaxJwG8OVa1c+CzIznpXbRKG3rLeXSHaJ7DX4CV8zcNiAGMHoITJ4yVnfX
37N/s2udF9mnW7DLc/qSTW7JKdQsWnYbRGapHRrrNU3klRHJqGvEIoW4zsPoaf2StK2zo4yrodCY
UC012IY9PiEdQ8DE0kJScZdHDSLOoQskbsJYBG8rLKOPi4IZTX+/CafGf7Ad+Nor2EyamnqZlXX4
8JSPUAufOdbSDC36rNz3PTyWfpgK1mSj46yMoy4CRibB3B3/Qmht+eqqSp6xaFqY0jogNZ4xP0Ue
3ediSXWQvd3GDTMlC706qezptmfnVSiK0KvFg7KdG9Q80CeglnuR0H7iV+IFWJaRZMHo5lguzHip
t0duFWQP4gu5p5OFbEjWq5KmtBneMqgCvwDBPl8ijRanbCmzYpvt74SqhXQE/FI6aOlBZZLuTHW/
FVrCe7RxT3AEPrnspgOBu7DfY3kUXleUMkQbQjjXh6wOyWiZ7aiIGOn1uaW1kXIxNMiHamJA8IM7
4KZgsvF9xkj/nzf5apzoRlWLqB8/NoSmZaP7fEk59Z0yCxE5GeqhbjiIWq4WLfqPDkhFbdU9+bKe
hLuOx9BH9rl15ycgcKKURh3hvBqO7YZYMj+hc87Pr4n6KfUmGed79vt4GQlHINAr5rLsOCHPJM6D
qLh6ni9eE+7I1zwqjYe2stAkAUwQlzfjbpP4D8MILFmJvIEtZFk/tXfn83x1XLhEZskP8HSwoO/b
nJ94ZmpEinFWcsKEVLuF54AMwQ6eRCBkeHLFg2od0rI/pNFy0EzzdtM667kCJrapN9aW/S/tDJ6I
43suDFe28NAfS4RziMwLI1rIsb3ctMhIYti8tXcvP/HbDVTcShcy/svhqmKOS2QIc7W1GJWa9sTU
1P9eokZBgOtSSC13WcIQkr1BiPtMNHW+7WOsDO/1orbg6YQwkUW57Q/cw747MmH5yZqKMGHog3FN
w8fdyfNJO2360UdgbU/+BqKfImeUiTdtEp+U1LT/tkRO6DwJyPgKj/hqVOmt1crmtXsmzOrfoB6I
OixsSo4p1KHdT096ekhYDPyDO3dA7UmE91hnNjN8ndkSeKhMwKNvAjMM1JixKcQpjmn/eIzOXeBj
tdgglv3HeYGLoo8G3hfKe/QUxHWuJVi3TIDucupoMfK+EIkty7nO8bedqzIUrBIVSDoj/zV6ulev
Tq6M+ACCysjptyzL4WFBONQfLB8hwj0Iw7IudsZr8ef+6z8o/ui+bWIRl7N+9ilazlL8xiV+ZVWQ
l6RtrFruopJri6itDCTFxP/qVzeOCfJo9PuWv02z7YiW4fPGqRQVcl+ITF1SsHEXyZACJs6pBJQL
sAtBIOT1XCAXPTNtwKAf6CUpVn7PLwbL5HZGGdxMI6X5z6fOgyokun68yRXI1fYJJ0ywam4GUgPd
+6bQKR5UiRRmPRceWoq/x8tIkwTYcOJ2BMT4M08SfmjvpHyRyMW70njecUfIMIar7T2yJBgVmuXM
HCnGyWyCEmICPQ1IXx5DlX8A3KBnZMfnRzU7JvQ2p4WsFhaOypNn/HXJIkDFu77PPFwG7RDJXpFW
RY9f2g0DEHqQ+XyFHH9mQs64Ca0+3mPT1vB7SFrDl5Y9l327Et9MGUfhjbx1IRhQuf1efXeJlgII
KNzDavUVSonzKMnTbuzQJNYIh/n9TVC0MSdriXNmWrBmkKeZeHhZekGyhpdfE251+MGrHbX78sPc
7QBe4fd6lZlc6SAbmpzv/QYtRajE8A9adCh9kcRS6mGRFgVyfV00YKSeKydTah2csO+/Sq5HJkgY
YPrKWcECSCz25rPpVVPQYQw0Br8cn6RTeWXatouWBFit8rz1PahNE+ee2H/MyQ1cW2duEVf6Ptyl
B1hzPY4ppSJRzLccZ/MxoPpKJnM0yXnb/6nWAvkQDHe3/qII4hr5f2ae0La5DnLkAVeRhoFnnlKw
Y+uXWxDrmIwhdA7HfLA90PFZBR89gmJqeA5Ir54fkwKAisu/HX8dWaXabnlbTQjHv6ak2UEmfyl7
xbfNhubbIGfPboHeWy3+kBJm8Ifehh+o29pfsfbwEwE64voHKsu8GvDMkDQExNCreQkB5snoELFH
TNBNN3Jz2hqyo9gieRdfZ+Oste1JlfhTSQp2qubjm2qfO7YboKEE065syjeQwnLZkZ1U+G+MLtmS
1u9z+wM4T2Ss02a8wN3z4+hhUMtFSD12vig0yF9+P4035XeVjJjIwc195P6thRtWU9NytB2E90Di
zw/EkK1P9qx1VbvO3TohXEfxD0sRgFnlq/EtdXpAnJr3cOLitXjNd//39mA0WUY8A9/a3WUHYOim
Lvt0wFX2C9NYzYVLBucxDSsPuLJT1Dz/yMCrrMYm8nQUGrQQqxzZwGwNspQmwHQqtlmzG8H3f2yP
YmanUNVhM35GulgNAJ6pls0ncGJMQPgSaqziJItvubf/wGW9w1j8wFYf6WZUdYS/eMCr0o41Mit/
S5ayFQ/BCB4nFjTEwsQf3USG3YDit/5Tt0ugF1PbW2QfskzP4ZslOwzEKdW/ANikX70efdJlUA8R
huptxRJOvJWKseaeU0kl/8CxASBDpQIxtjBqA/6F+ni3sr7XUtepBIDeFFgvTKfBT1EM0fobic8e
cw5+2LINZMh0SNRtmxwHwP55IdyI6B0xJ2sg02gnIncEZPjcatNuFb1wre+X68LBFAT6wsszBGI0
ntOxffFy0Lbe/knFtd4MOAgYAqwPIIb1R3bkTGGwB8SmEK+LgJ6T4cQilFjW1uuPfHi/HgyRCecK
R6ol/MG/Kon7Sr7RVwD38nOnaaMVsLW0RlkJ6RzJhQyy2wNWYl+Kw4O/+/ciXO/o8pCxYKK6b/gK
CLcDgMbz4LCkqRRUAWI+hB6sx+jbmjsW+NtAVkZ35D41448w978ohgEPjZ2gkAZBmaD68GVNBKOQ
r23sx5DxTG69wmzyEycx4tVIVk52A9ZWJhAtN/zyV7iGYeYjDLv0/hxTgt3jIThmech9kJR5BI04
hHZdyLb3NDp6otjpAqZzpTEvmQt0gtgXgrjTykhuYqZT7r8AIj5k5IwnGxHwypLpcKIj0k7h1zpw
bmwVrUd8Q45rP818hFWf6JRAEV8njVoBOFx5+azi94N7x3r6F/61LOPBAa0108fD2gY9C25wGir3
enUmnpkRWeBvmOpIsmjwHDhIUGfOzHS1wlHlndqDs6eB7C/+d1hQjWK+41zumCD7hF2ljgmNYxUU
1/JiTqpsazzmbyBM0y2/wd8hs6eVqXpUB07VxEqvlbKrqESAvVWtGFgzguv/ddU8GBeIlpCNWMdq
gZtSyOI4EgSebq6ORMCTyITEWYPEDBZZQRqXIkFMhLw5g6AkEW5Ms8rNlFZ9ekhABNqO0Ne0tJ/r
bGgpvNZCBEe/QzxaxZ+Xz0PAE/KTHWnHQOdlg6gl9qAG4VJ/jTNnPKYW+Ga0sVGrsjyGtkpZHoZA
39TE/UMiyYAAardIL2kBT2fw0P1z8hzXOSE2APTGauV2tuWWWjZ0c1HS0l/2n7ukegbZBW6NcXs0
I7NcMqqNhr1d4z8AyDVSrhgtNOQvxRK69/+aXto7Q1lPP3VotqPYGSGY3f/8LcaIwQ0Pl4kxBGTp
GBQhU3N7D2S5weEOwFv3+xF783F0AjO529k25/mZPIOokhJv2n0tTrvAUsmhZ6FtiQW0MKGqs3bR
LoripN4ZIuDsIJRwJHvfrsJ/hDMXJ78y66FMyZ3lxzTZvMb+jLG9789EfUkBwcv9omOgK0ZZGfgS
jtBRkdZPeVnKd1hFPgRXVzn7bXdssvblnSN5Tn1DLKXFTDlgd7NEZ52OuuvyWsoUWJKmV/dRHIUT
fPMcH5ll5lCizvZDpC92nSVOHHLCemCR2E4Yw2zl33BnYu6ZvLc0tIzhfdnoszhxB+ri7f10mRhT
AtnY+n6w979LR5bI5zSeH2kqfhXtTTAhY8vL23p1WjpN6Z50isqv9DL77TK2hN9h7TfcvbMiYwus
MDXQO+V5Bn1GOEk8hWxzG1cDST8Ozsv8KtyhAYBT6si7uE+INjb9nqXu4VE11xzKsmdfD+B7iPq1
L4lq/WOwIGMm/CoUlgt4xBk4cz+Z5XaEKemN2Pdr2BXsCYWbSyaIDJJn0qzR1vmnjtHLRQiiBsrH
RtunTjCPMuSYY75L6ksoVP4uPTeJB/kSskxzdYiMlmIguqdIPTt/S75SCkMl03NePhqLn4iWnAmE
cJFqFp4Y+KY+cncj7O6uNqQMQdVr94ysQ4SLTCAW00J6eh9vlFy2Up1mCG23ru7Z7XZdbVoRMN3P
qS4G2SGtWmDIm6Dft3qzi/Dz+KFoahibgTC7VdOtxekiAGir6XTxpvuaplWjk6kSjYP7/Gnaxo0L
xiwDO8SO4JXXYZAq6xoqct7ER8HqfW3L/EQSdwiQKwU04wxOuJPkhHMJb0Xrh0BMkF6ljCEZcSXX
jn1ZEe4ak4VbmMwIkNtgSA50sy9MhSin6CcgCJAe33end7Gu1XF9fMe9/2C0HlIejOu4WBGIgJyf
z7xxIhDjIQC5FIeUYtPC2IzzLKYkK+J74MAdVIRn8jIOs6wuebsJm59JN6IaD7wQ+NbYGnSbN8Oq
bxCHLBMn4EWja2Ff+OSG5Q9Duo4ky+6xKEY1sJEZdkG7xCpad7a38Lcwd1QQrWTJqSX/yqne/S9M
8iMzIdu45n2hzrtCFqZOlRW1o5qmlYRZhpt/FVqSf2VsHGJjj4CKTUGZ8oKaFh742MeTFbcQS8n2
M7OAglPDEuVw78cSIhuwLjRA6LR3VLUkr0dHfD+t6x1Fw/cvbCOVjuj95e5ZUp5q3ShO4+lcfUSE
jGL3WO/+RsHfR9nltn2FtTQBOoxDBM+EY4s4Fj3Ixn4PjgzKo02Gf7o8rVXnBqSNtcETNlCSxUYW
yG3iKYdzNvYbbtxbHFM3WpPN6HXDCQOzjchxkdhlv6BbA/Uuy7ip5EZzso5QC2YOTjaZx14XXIiq
h68RQA9sr15mIWEvsLn65I0fu5yAx5/mk/BH270Tlgm2WgoYImPFi5MH4nGMPG0E5axlDJnp8ai4
Ci/TXaum3hilSvs2I1SMmkSBpU7iC4SOwpAa3V5b23qT1J4XZebs99wb7wdmgwknn607oTBS4wiU
Eyfo9OiUrl1skhN5OXvKtBTVNwDSE+o7QEiA4grNksNPS8ab85IY09M5S6FpRnbgcpuAiS6FEh3z
bJHOGWDED1E7E1RC89qhZjf7W2ERLoC74IJhAk5GhDTw216Rdjy9CZvMUF+cwQaqIV3ajO4TpPOQ
M7mXSqszXCkzfpxZLN6TIjElaYiOmGqL8FIbEohfLK3Cq13MIqtnKmXyXLIJPLxjkhxuH8gcKouY
D3zkuFizp1M2w6VupySrATOzyaxlgnMjG7Dc/M1nlf38YBLLSllpxxGefBdVURXfvofVblvqqrZn
NvMvMSATNcH0YKZa5gbBGw0XrV3BkICtEGwPhDrpY2u4DUQBI8GAwlN0JDDN4qLyo73JyiRZKfKm
ZelycnWHI+CfYJe/OcQWt8T/EsELjdl8jvdgmXUF5mEUlpk8Sp88KSpoZZNQp1ikeSaBUPAkrKQo
aJVGHuLs/ojhvo83sAEJKYTOTksiU8B+MC3srbi5vmrubjNlShoJl5DnOdFb0PNKQz+NHFAnz41b
CGDBhOlSMCOi0aUZPmxzvfkgY8/+hW82DCk8xC49eMcK/0zZV9YFqASGKGtlFOGlDboLNwB3rHtu
lhliyEtWrX/3/x2JnuFYMFHZ08Tj/TEF+j7zlFn4NymNxTteLPOhT/tPHc8ZNp/YXgyOfklXF7Pp
2p9+K6pzTTdKMT4UEz/tNR6TSxc3dZgPqGWNADdvfcEEeCGQyRPDGbqElGcVAuo4q+0njCVrGRvi
4KKlgCUhVRy9OZK2bMq9aD+gsRsQYdFj6MeYC6HUGmiDYlyy5snYNmSRgMwYqDhmJ1QLcL268hon
n2w1J2iUrT7BmGUUpxj1sTIEJl4cXUs3T3dW6irQdeB+TCksKR7dconW8sW2IRTWl4xhZU9lM/7v
PZx1xxUSyzrq3UXe6Bev5QCwOxvSLfQ8EQZr6SlaVcYQKwxxn8m5/Y+KcpkNykaJjBu4clTwEqp3
hrn7vidhjwylmrOrUFqZvzRDTFhdl4rSD9MrLgbgIXAPq95uA9BBYijsiqPPwqdy9lAOH5H9XEtZ
yfLpjznyFYGTPz7fmocWjCDN5Z8zXSaxr14nqGlUKMq+TcwOlFxM8XAY8ITFgnOMP9/uo+fkBPGB
T2n50eLSuv2+A433qAG6SLoDXuvCSFG7q9RvPmlpNOnal8KibqwDwRbHvjyuRz7oT1ZeKhIb5pwP
FTxNpXdjjOgbbnaKH+OLzOSJ/cTZoQR7NucQIf7o9xlFXjquH3xODHZ6Hr/0hy0Lc+PZ6JiNf5tZ
MTpzseWNHfJ1k2sUJcZtWZT6fU70hGOtPJyKXb6ogS9rdsGAEy0Gm1tPM09VHyvMsPjA1jrnp4iZ
prmqYmOiRDtjkfVsEPalDfHdTYnNpGy8UKcBuPNGj3+OHWChp6OCPRnP2BfDUQpR51kz0vh3XHJe
TUBE3ONFRP4OVbBj8LDIV3xv+XhQ+L1t4vr4NJHn6K959oA0ZGJmumILFK8iU9yC5Oz+VwaUiZRJ
SEpQ83Lehb3+MvD1Iq+I8a3cLAK08/xykVz4mpdymBsmWyu24a4sXbgxcsA0P/0Ekx8a9jD8Q7lq
ddIMHj2rPm3ENEuDUgcZ3m8FqmwM5rkVGRaN3VM3q7eeuwOkMbdlowtV2WhjF1oCbIxvHM7E55I/
YdGYvn5xBFeEdZR3M5HDKiDA4exJxcY0loI8ixU0Tt9lxsJIn8w5dgzmbx2WGNTnaT5cutl8qO64
bns/R+WHNOdh1V9aQiKH3tGFTlvYdy6GafL1ZlshcE8hhr97sYPo1SE5vhDmzoOFs+5ArnRcf4ma
6cirmCekW6oLk5Y8w3HATsERYUsPsCHtUH0AG9j2rvF/iVaP6l8uEvxSQXJYNzHCqdp1agmS8lyW
wEE+7NMFVSurC9kZr2gFSGXymUBlb6Z9x+0q0SW/Tnxk5UivuY2GVq3jl6r65f2UAGjjgDWK3/B/
mI4aw3PlrUz4x+cLmGY9ILO9sA6v5BVtYBNRCsfd1A4te2IgyZNoVUf8rmejmagf2U74Lmw8cq8r
S/Gg0XQqhoBobU/CSU4O51Oy/1QsoDSZ9hGg1qSp9dv0WdtrJSZJQKvWxbn3iVOHA1mqsqHLuWu6
Ni415nioHsxrnvrvBHu6V2prLGi2ZM5bblUyCf0cAj0F9n4Aq5XScH3xWBiO7YPrNMhda9UVGzdI
TbcYmmxMpK/sjGqScKwrhfBOEUxTftebvwlntzsAffkoJ6KTR7DPG41R0CirR+qiZ7V6dnZTWBuU
vqMGRJKzX08i4LWKEJ63n12VFQYHj+kk9DHgEiXRNqglyBMrC5IilF3jk1mJNcHUtBjM1zvRCGwT
Sdd5rs6PC/EQpRMuPrcOw5mXxS9AJdSDP+KArdCXErg5eNGoRFaauH3841uw3cnvxL+LmbqjhoZv
ChY1AD55HIhexte1eoRUC2FWbs6nohqUV5Dsch3IaupjlaTwAAn16VFKjBF6/9QMQ1atvMaMLA4t
VNQBvQxuGrosM1QhcsOlY9XydR8hPRthjSFlaDiGlVe1S2PjD6RtkeLWxrVNAHwEouTze7EHYlds
zPhSDfrpKoYiq11Xg7xuMlFntbypnWX1uaTWFPrdaf8e0X02c4mMflQLevqzOs9FHuTzsrhneFff
bfYAsID5RTJUinVxjGBoM592U317oJFgBNCM6yWB8nm8maUbSOwruyRMjx/YKeEt34prXPXSgHvz
LVdppyz8gBSdTkbJ4E7i+HaadH1w7xlLOJOacFbGQ3Pli+zmmDsHAq5D6kla1clT97gCiVMRPmf6
mZBAWwGisl5DsafQk5AkUlwfrt+nktgNaKJPQ/k8XW8Hynawp4M703uZrG5h7nI3pSSdZEAkCzS/
trN3JuKg30v3FRX/+lveKLC5i2wEbUCx/Ez3/WgIW7DB1j0dqRIsxPsSZcI2JXufyW8weECCBNOO
64KnyNmb3zn9kottCGgNEVt/uy9Kedr962oRaeU2uGDxb2d2k3wmH95r4ZLDlAG0inQvCA+YvWNH
BotJzbo3doyaR69/Mbs0AObLdgiA9MmiTMtf8I3+3cyfV3GM+b3akDAleDnrpql79pJeOZY72N+s
xBWHz8TlaPMUFtUurJQTIHtaOvmmH1HuUKmRwkBz0ThzldzH9q1XyifF1sO5EEm6m5531ZloTSJ6
VtOlXSfje31TK5U+9BN4v5XIFm6QIFUAdaEUp1RixaWNVQDZLSj0sDV17vqrKRwkyvebAYQwe4QV
qas611mZnUEI6X5VSmLtOJP90X09bEIoix9bqNsyOKZ+8p/Lv7JgFMQEGGUC6Zn2SVYhrMHm1ytE
J/XDE285CZuj8wbEEEeH3LLichR87z4B832eXAyslDvDTSMX0iQf6xWiegwh/xnT3Iw1lKtJqIKK
3mU8DYw5cTdXFsyTi4ufzNjjXQHKfy8LbEcJfRa5u3hJ3TbKP9hI7xp+6VBfeh4be5HOXdNan2om
3I4Ca6e8xkEHuLEaqK2kWtOkDJ38yQm1EfT7qNH1Wh316KFA0yTJXqsB/Xo/FyxXhrU0webY0/am
6PpfeGcN/qiUrqZ6/WY4+rqQ5BH/ekfRxtLJclLsxMqyaT9gWq5F3Oq1QCN8Wn50ST7k7JyH9B9s
ecSx/KqLZZbti6vyGdEyOrdeTBJA8T/BwOkGRUKdiHP8g1jwEkkUKUqNEx42RSsfMUQhOb9gmt9n
tDIxynzp60h0AZf4pTrqckR0pPUJLFc2YKiv+j4HUpzR7l9pxu7gHP9zyX6ITLU2dKt8t/s30V8Y
wzP+0c5OKZSDqPlbl0ZPMjilvVzU1qUO1MHuJW1ZTOV5POllSUSBHXBeZx3GCOeEqIDaXXfaegjh
BusdCKeKEXfjxmgqrudHKcCyIwoJyjzHSoJ1wyQ+F4FcSIKZaLhI4uDz70AXU/I/eA68jnTsiEgk
8Gl8Z48ysFau+UPzJI8H4+No/g0/eExa/v0Ot3jHZU54JmCxlY+Od3fYrTb+XwnKbITk6pMYmeVo
TufFFDkyybZ4Qkea/YrHHmh1Tu+H3wHhMeMXHCOr2J2vV0bQYlYFbBJo/UCEbp50bWVT/AZB1WtW
1gR/FoeMxo81oh9DK1JhVjOs0dFybVoU/dLmPj1CZp/+zpQMdPvnbzIgHaVkfLVFynpH9bJRxlO7
6/sXiD0sPZQXD/IMFhP74XnH+oPH7vO3Pk1/06k6aqqS5eiY30bAQP2Ah3GIQojuFeVTj/00wx85
LApBBFEORRYrYXpV+cPKfhBLN4UFDVCizCYJFrXFehMKufiSVkslCRClpH9ZJi6R91YA266hWRgK
ggsQwu2lBLsdvSyxQG0gfkfk5c7zzyt+4PQ8riphC0Y229IjMewn2mFy/ZS7LtOf07QQO+WW80E8
tBHlggKMSjeYDf19dopBolkqNj7GsdZ+qQuqJTEzWzKhPfSIrhanZXTPSQujlL8fGvrYVY2Y3zcE
xIK8F7v4KAy4fV0lZz6BTmLl696KjN1MS7X1w+Kpg7BcXSXEyxuP/Ms21vtkdS6SP0ZHdMmzHm/l
C2d5kmDJKEMgu34TiCxarMqEzUXQfa6uECxLi8zXrqW66sRdEKvxB5UP6mbZbU/D1ZhGtp2qAgC7
Nao1GIV5lfqtNAr+hfdkNnB27O0JlRPJi+SKmFrrZEosbVgjzIQIidcC7tJZTqjjPZzTwSCDHkYy
SxBz1R11Yqmj+K1W2TWF+asqNvpGmFMRNjsc3j7kvUpu1zmaHwb9vWldlI1Id7Pp7w21GOETfz62
2DGeHHOqJOC1DBUwywbpRbV/6e4AnJ9KIrUyD4FeDpNQkGPPaL7qiOXSX994tmbtOd4kctDLfTsV
3ZGPgvhkvQ3UWLi8VaJ7jlRAub6MxYvfn3v8U1IBp7gW/Xo8ole+lPDArThyWfRz2M+Guuc0bbQW
0Ut8EGHfDLQM+YeeKokVCRSij7judAHsbV0HNIx9ERHYkPqhiR965xk2iza2f/6t3+IA2fWlYCuP
Os454wXJEuMcVKEBH/TezQDStsUHflYU++Y9UE/SyPkM0bULcGOAlbcxzyzXuYzEhoZs2L2Qxmec
5V0toH5PibJTy2RJfY/2nA0KqMPkZ5vx/R0BwcvMgkTgXpACOQ1yc3z+j7M5uX4HaRKuEswUbJ2l
YpapJBVpoK20mYJgAtKYsXWyYcIc8sBs6IzL6Th52ooO3Ejnj7i/85y1Tuh9DsuriQVa6n4ZEbAf
uAFnGqKRNJNR4PJvyW3l8oa0fmhMk6BnO3GOVWvLgCJZwaanNs+bndr1ZUgg+Z2ELwHrkGo5DUJy
XBok4m4zTEoZXivQUa0fjC0o3JNtuU6TMLVkf4jiVqxFb2MbATAenlRH6iESE3U1WfOJ6ksVA0HQ
KkImAjSrOTrYMI5kIc6nZhk+h6AU667OlYPHixyStwJ7i9B2gtDP5YBcKJQD6LqKUXqM3F0848ki
9NTq8EW8t2C7aegeTIKqLryaXOsr3n8AZpJ3Vq/R0VFh+CbzADf3YpPf8rG1Arij1MBwgiCxtkvj
qhy/r2ixJf/sa3+ncLe8GWR9xakbcyzJ0V5t4HYf81p1CZH1/B6K+BBfFhCsiBbWWi3yW6pCJ4Ec
fKWqa2PWMithuWJFg7oX1bu51p1RAEMarIJ2ZmVDUMoOa79wQKPw/h1kR9Wz5GUTDPWYuoBwgtm+
NbWVLAhSRIHw02nWE+Ou+/GmNI3Cuc85HWJodsVQ9S5Pi3EwWer+CpyQpiGbYTfhjGMQZnPYBQIL
2R+LoH0FDGkcuSUTq5i41lvPcTy/KiOMY2VQ4jV1BZxE4PHZqjoo/zgLHOYeWGqGHtfu0VsYbljQ
7+R6ZFwMaVrxADM8ms2v6r48QhD22hygttMQaGPu2+v3AyFZ1CMxHJacZXtRBJlzGiECIQqJiJyo
IC85z93ptGI0tc69CoOeDodH4j41ooDM8fg4JacrCRdOk+Z5XYVLF0uuWSmmXasd2KeBnZLjkc6B
dDHWSLpg/JXmvM43r5CXAEtXdeJet3LV3I00cRXUEzGn9jq/UbipIbi1wH/LMoeFMgSl8nSv6iy9
DPd2n35F+1dT6qawtlbZiIfbc027UXktg8RkbuPHI3YmrXJOswrZuWghIG2kT7j5YHn4olBZKEQh
K/Wzxv3MF4+tyCsHUNoJ+YfdzFCDLn4YJVe6R94bDU/OEtE1juq1BknUcucV8mQs5yNrKySQZVsS
ckiSxWGQ3l8wfy5isr1DYKPWFbGyjtXKUygv7o9l1zSepCZ15/82vXrCwlJtqdxKeg1Zhr7sLm4B
KoF0LL+9hbw4QkLPQAecQPD0smKIlfHCQUG8B28ry10WAws+CBKA3WmTt6X3xmcekNPqAj+5fBye
+OsJQ6E8+AsLOPRi1FwCZoy8WTUIVyXS34m/EsESsKtu0jEZTF/K8SKgm44syvhzwYUYcp5aBrHo
VtP8lxEcF2Gm9wYlz4Dk3U3Q/m9kDdc03F4W+3h2J38O1cctQ5SoEgF5It0KWbJs8DH8qaefPq2X
xo8JBHhiWyZneFg0DJKg9ANJkzrArRUWvvYUegqb2PxnT8geCdDN7+vA+mDrCKXND+HAlGQyf4ad
u9hm7s+/u7ZVlVJeEzxYwux6oBdhe7NlasnyY94X3ilzUKLQqogReZKtZJHZdY7Gt59h20NtlqJE
Rioy1dw5d0e7SMH1A3nDHTXHGal822rjkjMf5qMuYr8m0vPbPgcuG7RklJzR4N8/dgKWQRGirTWP
sJlv2DmIiOxPRuLGMqX3Icu3JAwS7iRFz2oYKtLS4blukdeY2jH2fYlCMrsHL/OPIOF4S1be9ThS
bWHkQZCPO75qUi/+WlJE8r05f2dNRwGnWWKbs8+RcR6e066SlPVi2aw60fAbhi8Oxg+xXsjwl2BK
FnbfwV0LoCn8NdcwCInS+EF2eYJN1mxaqZDtOeOw4TbdG09/abuFCti5XdtglXEEjkzaJfmi6/jX
UmTZQTc6sHqrsrecjziEppSViEQv8XIhz50AT3pJP+UZrYx1GxTKASesvUwFxiEq3U9Z//i1mqJz
+UlEn2xJBSGdwqjYob/rBFqXJOgptNUbDVE0MCkD6mOb3r7/nfeKmwim0abn2CzErMS4CCoqors5
wLtiOdOlwLf8JRGsfht7xwJT0F61wctCYMi5LMwh9XMC8qLHBA/I9lA841/CKEig1R2NfFdB/g52
pBT6Ebowt2rVyVEk/0nBUdYtqDshenOmiadhJvTfANX0ffXsvb66GRsYlhmUvHurFLiF2QaJsbN3
uuwr9d7g11nVvqhldeslIiV8mfE2/t9K499d6cBREHAvYZISF9j9WZYNGiWZQwt/0oOU+pRFZ5tn
4cU2YUAQzEioEH0+pt80Wh9UkSHY50HkcrM1ESOc6AyYHR4WUuQUcQmoyAyT3s144DDpeg2o1Vql
Blm+UEGBfdkVsNnHXy4yFRLLmpng7K59OKsg/SQtofK2JhJL/fvOdeqtqLEOmpXJEPmYI6L+6WVr
ASSVub49k0kiBu/vUXTJ2ZEj+T/7uVP1Vexu2NKOpSSaJVssNZz913/qh5ADp8pxqTD75XRo75wi
DbdvaAvipBn6TedZAc+R7gzHQXAPoVeTAFujZycKyjt/85IUBi2bwU1xC350Pc3cdQAgeKKhRIx0
YVjU/Soj3uIRBz/rQvS2kqBy0Rdp3x5/WS82IwIVLOTdXIwP453Y3wIPE4IO04MZ7zUQP10JjcJj
e6PkFzj+oycQDRYYbfhSGttCnq6+Ng6bT1BvMxvFDjPsF1tYWOUsImJXmPdaGLmaW6juOmdv7BmR
8sKDch5jJwrLxnPHxAVNbilSdWFuDR0d+G7QzN1ueuFb+xT+aH8cjxaz+dtC98mqhUIfVK0VY373
k7qTqwxyoZyWP3IgbPYhe+XHXVA48zuPjXwXbOBRDEHibuD464GSTjKWHOUFEzTJYwSU/0NPIxVV
b/mWDT4sBMvbRxAzUMrEA8Uu8B8PcWmc/Fgd66kwgr2DC3xaFOzn/v2FinvK4kkwjK/7xKi80ZdH
hDBBt+p9eArVhdLAkTNznFooLuqEkzNkxxsajRVpG0xeuznQ4TTVLHXb65RfHS9aIcm8Qxt84mO5
Wk/H77ZEloxhf/B5pnKrKpyHMrN7Mlhh+PRaMJ6jRmyO//5vHD2vwT5LE5HjOdDpzbiY5/QPREeO
YlhnVIEXJyIVOZGQZsz9jkqszG4I3ygQ0cp4Mc7lQ98aZpbB3/zgQTcuxL61shEDKOr3grGOKZFS
6Vzmpi6ypqfPuBXuayoD/JhPbcbt0WefNVOFbm4tFKB91Fo2mxA6jkIvzltIgcOuDkxJo4nvf7Uo
7JFqGgH+whbvBis+XpDw5gXbmzxW/yovKJZ2Jdzsn10c/6N62BPO7vDASeCARegg5zO/IMtGFvWs
RdbSP44iECHZ90dPP/2sb63D+9JQljLp3doxkqad+8A44cy7ilcctaUalbnNR9rI5g4RyrD8sX+7
6YqJlpNBif7sDUMgCwB+95D/KL7CzScwUh4xhPtRPcVNIYQiTCKn0Occ9IL5PK0Tck5aZ2DJoZIr
9jrHJ3GicYdiQrUTHz0bEg2XYi5HD+ZN2qc4HR5GhIdYrHw189sHDEJzdDOj3jeNbNA2K8dgmH8k
wsNBWuGQYhzdBtS3rUiGX1F/T7/s9JiYpZLz00DPNHsLGt9wGoNuC6kIFv2y6Me2nptf6LrX2IvE
R3EW1POauMoqfGvcJI+cLWt6AWZ3g9wTWhhrja9/uQKgtXGzmV/JOg7j5lSNZ3/YeiSLxhGtwXNc
+AY1uxAcLdJhPW0KEuu9Dr4tYtM/2cTY1LeComFyyLne4Ll3upWzyZMNcQFrbx8T2VZXI3Ob1DuA
sv76UwrzLrkzSg4uR6UqPItZUotMwb/C4ChrI02OfnxfVwjUzHWIaa4tp7BKu7gCY4Rw9AP3hRlR
cckm3zIbHNv7OOXfXpaogzKPjHlf2q4PLsjfFCpxDI7S9iI2fMUr7wahqAU/QHpDMPKnIhYqwLd/
taociGGDQfafbaSjOOjCX1LWVnASJi+gTK6B2HAu14+RCXH8PLa6sX+lVrNrmMcR6hkDjTX4WKsK
/DXC7jcUflsckNO3T+FddMC7VV5RX1fvlfZYacuvrKT16sdDtO3UTGUi6ujvTWHYQwLaVxA0WIPf
vRaxQ9u1i3j12WUZT85OtM+MmQsVIma1wAnnfNGZjEbPKkOJ1JEKO8TfwGsArA7diQ6q4TLCZGqK
TXez19nDz4vw0FESmHp09EHWsvAFbIe9Ws7ml9sMT9zFW/TdMd/mdPQcnp3IP8fWy3/SXsYFOPiQ
BcqJld5sWnbLm8nuqdAY4GgInRk7Ue6miUIXQTPvHCNtCU6O/1f7zJmt+rMsDxGSEZsKGzksah8P
Ej7zlWTXyKTcegiMMv7uu5Mwy41dxh4O7Bv4OAIvGljmYxwPWAeNnk/u18Mn1umN54fiVAVsDtYe
8sQmEzXQ5+vSujSgUnFpZBJu8wNNXO3GFlsIQcLYVEVMQSoHf9jVc2QRobt8HztL68FfhXOSM4/I
i53mxowKZZHiJj3TG68+GVzwcYhPcie64HCE7GE2Lb3K2ylovlX7uK8wJc0v1l2R20rpDykAxWOO
OpdkpDL8MTWC+WQdbwwGYaykUOoTesY/sMirpB5tyqOlQucm0BKjoRJtCR4Nxcwp0VfGrwXw0l8K
lpG3FAfsunbOnfJFvylOpcavY4xSBijfvieSdnZPxRjwozGb1CqVlyz6nfSZI+KNwkttrLMQUw8P
cZifzCMX1LwXdN5LKwAlLRUYIti3dCYebU6uw1piTGiY8+XYuBnO+YXvM1aaqtGRt3VEvhws0Blq
+LZj5VcXUc78dWSgbaNH2ncaidqj3yzjJXJArc/MHJb/E4BDXJdCbg/hogK36dppSYI/5xB7n7YD
r7aaa34K9QKCuQ8qs00YkXviaiJor4Xj+1gYoi3KHO+vQ7TkUBjk8dEF0VUngPUW/hyoK4F1Ybgb
MunRLxoGUx+KXOgb/52CR0++4kTzDteHCmHnlx1OUbIG8wQw+E3XS3IcHxRzaEAJ6KraMTEhIOR6
e5xbx3sR0Bh4fof6EwYC384Rq/XzSefDvVlpg9+hBX4gl/OY/yyJKoWkD/jy3jvYqXmhClR6Mzeg
ZXNf/emnlpFfphklSAR8quWjQR6mSEnN2nin+oJxBTD4aAa1tV2oW9m92YZhx2e2DA4Cq5D5OEjA
U9wlJPCE0IWX40arV5npFZHzPki5riz7+Rc9O4tM6AeNbjZ1Pp8VTJ7EiwWPdAYWKVYjXxzzPTmK
kTFd77pDjlrFrdiojFwiZQlXW6Y1Ra08PD8LFS+rS/Ssb64KxJQPT2I/CwkVLFUs3DpVPA6AFhAp
aJWmE4f0VvcHSEFlZVnwFBJHVSUTyaZ/AQDcsHmS1Cx+kgFiQ485MbrJ59sVHtkz7OCdg7HCN/pS
JWVVhXmBZx17RTTSD83DLRYzzXvXuSRjz+d1zurqS71xTdb0AnBYHUoWNIgqN27Ax+xFjf0wpUwu
Mkhum1Ftir5YG+R7e2CiP2drKfcLDOlOrvLqMqZEQd3XDjOE2nrHI+5TJi7nPGPTWUY4l7DQ9drF
8gD5aLf9FTa5E8gVwb8I/H9jmXvcW4S3mUTfuOs72TJY5w0/GunGLc+MlT74dHjnOsprNcYknbre
TPddWp+sSAN3DQmgD5tqbpB2TYAdqXGpp/7BfxiggN1soQsP+Wcow4wZ+vwbeUUNP7k3bx+dibNd
9hTGMZCq/lTCNg81vMET27rrYBEDz6MqEOhYKgLD1Jdpmq4vRCs5UpgmOU/hMovAvG8S8AlmBK4n
P4D9HXF8ysVkwcPOtLPAO04PnGxQ0SNjRf8I348sFlOkd4Ry87M9VII5PCvQG7DmQmgf/428in8B
S7VNJAi4dEaISozaghS21jkMKdKBFdkNi8BrX+OPPG12MyydpXzbm33kJKLMKZJeL0AJXPskMY/5
vc6Cgh9m/4r9pi8Nb4btPwEfrAJGOC5GWB4zy08cuyBb56X/HE3xOLrf2H9/QP8jnqbGhWImQQoz
37CiTQ0vm377yeWXTEk9ORLiKlY3zZ760Rv6hafaHfdXQNA+PtE0/fRH8yhxnviFD2IrOXS2trGz
mv1NsFKBOAaWXweR72nXbMqzVItX3h+IghovkIRlASgGfsQyrE/O98CHb+gjUk4oaRx+DbNtPXje
RW2Ychb6z6NoCd3otNkDa+zUPj4E1fgrnh4Awu6C00Ue5ezvv0v9mCdgk81dEYhLj1DHmK4XpGDv
OV77/l1xeLpXhKdBIgx1Il+ZB9Z84SXXK5VgYBGI4S3oBv5qOKvRWs4fhGH5JIEumYJ8OIgRJfvn
gphvNLztdFOm7JjSFS/WyXSqswwmxiW2Lf+melj3IUFZKh74aoDouoJgTeGDM5be3zG9pOsopFhz
VvXuw22LWmn4ClcqQA/6+HJ7KpESlg+aCJjRhGk6gNETgFwoIATlgcDQbwdlyGdUnM/WKsEz6Ph0
c772Br8+qI0WECfSAraeBD0r7NnPVI6Dxx9PhbwTfT/CqveSKoY74nL3iwgFDVPb1SF47zw6XBd2
DIHwpx4ZsPkuXS9zZde8P2TjJc201qNS9UDFYjIcGDdzACt/7DwRzQu4xm4kIF3JC5VgaBae2/U3
KHMA6K2VWZG5cIKkM56/cZAMSKa96Hz1X3EruKyp2GmkO7iD8wzQd597Lmo4kBscbcrhm90635Cz
in7fGSsJWcjxkqiG2rCCSGZo2C6ZxzrSoY61yZDut32ZqBhVaYeLGwK0Tcm+qjzfV+pMqyeC6FzZ
WyF9wOmMMbneDLRIXMzsIry52AyTZtSF/xikc4f+dQYTzLf4Z9Xwj1/YOo3VIUW8pc/Pjh7iSAqH
+qPiADSKkFLQCm7ktCKNZ7giFXKN7aG7Xp0adQNLhAZBapo7GHdFjNsIPy2nxnFUOwYFtyzfw149
XkFLFaI6yLMTB3COZle8J0fiqaEbn+fgSpRPeeW6eNB8J2gI2HkP/m3dWtkHhvW9Fe+wElFo9mRx
vdR4BmZGgBdRkGcj0mH8juZ7TpFteoNNyfdruZrHlYE+5drgKEoWHroDKi9gW8k/fVboKHYS7pjH
0Zt/j+sfs88JHyOfdQW8YSLmgHtQ99U2i4FkH+gglNM5sU2G58zF982YpXN34DhS+uKjYOJGs/TZ
UnuEHAUX4opn5FZ3kYOHLXU9T+uD0kE/6aX+Cz46br69mOgMKQtwCD6JVunAS77VEwl1TBEu3lo7
Xxmb+glHLoDboPgCHwks1XobeG845wyeaonzjStKdzTe0wYR1Dqp9Ql30/U1z241SoXVhyzZ9e0o
KQpaBASrNlgIxn5zo2kmKy3bsdLA+mPjz2glfBkAYQhi9W2z58iri9KowwxfNojcyXE+PbbHvx5g
/oUcUtAfq+gZbGE/OBiNtU8dwfcjS1G9D/yowqjLhTJsj5j4Jkqm2xp+BqnN/Olv2zCCWAL9nRpL
wznzRXMrofPMZTaw32eiJtBcBehxsdmLoeOyH1zw2eE7yBUN0asPQCa7zKxuL8vrxFrPb3AbLnYU
4YPWpoz4rAcHLMYkw8wAupi8yoGw/1S+dOYzucIy2+kE3++BMDuSilqU3AcvMmQ/ZeNFUDIGmSkw
TLMiDkyMV0VzsjPdbRgVJz/it3PRWN7qWSdBaUMDc3/QqYwd+0NJVcsy0aViud+WgzxBMVIBFrj1
k+jw91Sl1WNEUNxtwImsvRZZ0KZopqpR+x4Qa0txVXodqyUuZXSl3aEz6fVs4xnE/fe2DXNskFTA
4fN3tRyP4oVak5QKxe8u0MIKSxOXkJM9I+Sijof+w64arE5ECXyrI9gwIjp2IQnWv168kS42UJZU
08TBOuTDJUq4MCcYeSsiL33X70KsKiUVqPIzHzczv2HidxSgFv5f1Cye5ea5rTARZ9lqhTIbSO8d
J73Xc1E1qy5+qQMGI5X8aLlFr4+UrNOLW5x7DJjaXc8lFc7bpJlI1HWgKGL2D/LlbpAz6rou8L0A
Hdv8sEb0mkTlVE2XHP1QyHpudZdfidOq71UPGQBJ4urG3IZzxPFI8y6X67oXcHciq4OJrXAcCrtH
GGN/lTmiPGSGXlcqKmRbuV9N+zuqQXqKPjqxxsLls0u7Jn+5fVTBV3whAsWxtiX5Y56zhI6ltIgg
hp9pT5v8AJzIfV6VInJxHAzErTHLHtFjEbJVHvSuZ5xFbGTSIYkzn5eR9un41Dum3YE1Fbbm5fL1
Su3m8cjihCM/qVGgMhEVsV7FIkTm/+ym74EGEg3n7csCKwK26KRiYV8CRM/IbyXKlfoAVTGfkKOn
lEXLy10z89536PUvBlqMQk3JD/wbh3lGyoGXKxtQR04eOGaWL04PxY+8b4+9FyTDWq2JCfFVp0Sq
/6TdgQjsgA0MKT2Cn5TtrVuFde1CooCIXrBpqwNPaEiOQyaqISRaj6+9rSr2Dr/GC6Sh6FL0Vabq
/0jcWrNc9O/n8be+dXrYZm1rElmIMkZe2XLf3TOoWhvivHc43paQDGK6/YkmUlRooRImx+bGVueP
sauBx+9jt59owQttT7S93UbpJXrj7NvaIZyGLak9+6OUpJ2Zv78MM1OVVLGKPyrRQdtTbPMOnrHq
P04HSn3H4EQVqqe7VetDq92dtSqoMzf9jhbrNpTYaRJc/arpcYscOaYHUiprlgKqnQ1o8T45y4Zs
iKkbPU0LTnwc3KPJJVlmj+m7A7h25nNNvPkb7I2yxTjpVCygRfAhG4SxpKKRZJxRUW0keGfOlVtx
fU3TsZiZq5Bg5W4fsGZX5OpB/P0MMEvTvSoi3F6aG1i82A0w/DqswRjwzsAPcQs213KS0xbPoSA2
KP8XQWaVKTg2IL2yuqRchOw+wMs+ivkydKq2MgIXD5eBYLuZayXLOsCsBXOU0MWOhuqcs4/iry2N
YGbN6WIie2Rb5IVM8DW4/gSwWNwUr2Y8D6X7yhA0dPbTwgOpa4HoRGOvZ4IRyg3ADpz9ARcURj/n
D1Va/G/VOe7fVqBKyke8F2JgKsSCi7XUNGX0JzAo+ShNWQXPPF1TR2CdoEur+YjMjMoBhbJ2VNrp
iyZalXIKWn/Y3jqZ9MP0c5XFjwO9pf/GKeanlPobeAiP6yE4XAmFQFERXRuRf7iGe64lq6Mj7D43
BeO/73BfT8l/xjWYWKkQgJpeMdeATUkFbKcYVZaNO/++DxzszenqfFdRke1GN1HMdavEGzy5n6zn
wFH+E9aZ27R36c7SXmFX4NtE8yzIiSHeIDAm9dxV9hYUMrJXfgT3RGZfjPbYpjSYvcCz/bOHdLQy
o5nJO23Hejk+nQJrciTooSYFPXb7sfgLt46B+pxIezWxBYo3PaHkbj0/U46dA/00rqC6QshTC/+k
ohuwtIKerTtO1vrsOl5bfAEMkQ6yfaSk0EWO0zk5xbUYGfSazhMjbCw7DOZ+k5I5UKF3NNtDs+os
fgmV73TY20aszCFeyQNiQX2VzqNP7xRlq6fXabYRx3h3fRpgjP1jcF+keYrljsvT6ol8yZH9YRH/
a07Qh0XE9Pzez6E1dgUst+iD2qu1NkYIf1XyP3W/GSiNeHNEMp17X8yzv3XYYsGcnTqU0Rtwc3OV
Y4vjpEP5uvY0o8REJl1JRnpql/Tt0ghWtyvBGmZ9AmZluEQQXtKt3l0tpgtGkf+0FzRyNT/HoGg7
kpCPoHdDm/pbcgiqpzm7MpZ9p1bzRydlzVPgvZCdxcIzRajubDlgy45NgoZ+75+moAcgRJx8x3g2
YeRmrHQgEN8orpLASVj0rk5ZWh00oS6/fs+/Ql8Ti8E1SCDzh6px6e9SUUgJlg0yH1BrArjVZAEo
Mb9up4zz7qoCdlv0WqOBF+FDz/YnlibNu5rC1WIVyDV5Yez62QPexeJhqyD4OrZrUBdCpbM3sVVo
lmrI4cXTvCiFRJjXmBTNMUd6bEH+T2qWwUuNsXGdH7qY9cS/FgVs4NnCXp08RF8M8DUmgT6a2d59
pJsmT7gnhABZtVGNaSTmO7KyuP2Km2LvuBV9HbET6Fv6x0vICet/CiBUmFOpc+778xzpitn53bRr
wByO6DY5ENW+30/QIzNAJyZMBmVePrkTzKwPwC0nySQTIq1vP8LMjipqIrt8vX7ZjJqhKbTRH8et
ISwAkqpyEt++TYuO6SXzPGEzPmGbUhB5kZJ4OnmjfuXTo151+K9BS/KGGAl/ghNjQonhNIL2OzTh
odjNFYhgEE8gT0fZZNlmaQpUOzGy00h/CzKDAgPqZb8P0WidGVz2er5xK8R22sLWrHZl6jtOGsWA
bF8fROX+0F+ft/GfcFhi/rqojTwfOrO8VD+hllZPTIHFPH2ZtI2xmmXAZrTRbMpW8OXA6uRcp5N6
ZGCXrjl45TnUmV4CAuPVIrjMMDrsG/4KUB3w1U3geG+T/yLgLUSEBpBjGvmmVGaevshZeRptrPrD
TM/lrnLz0ZJz3fzSNxxv+3TN7yJTAEGBUMrc/ofBfIZB8DHyx+VKnOkOvZhMWjewHBYVCgWxPKhz
ZZWoh0zLB8ZYI9Nf3dZScgloqMSulvEQrfJFJfzMYySSwUhD4T4xh6qS66dw9zIluGH55E/d3EI0
V7Oa+SDzZcmQmoILu7It+pcmKXlFdpY6Olro3HtsGA+1SGCv66e9XeoL5FwrZCLGAvlJfsQczKY/
66bRC27x44/vgUM3bnnsStKINM7AQcXpy+0su4lRzLMS1T2F302qnpONg2K/bNhaiex3Y7usX8eL
bnYE/PeQV3xiAR8FjOz2w4J2TKMmjnwmaqIdkUbcIx4koe/m6jDt+JJCs8tZNc8eIFrkpd3b70zj
1bKVhneeHUWoKvBxkaqDzycdlpreH2pjyk1i53OsgVEyzN76xE7c5ZIznQhiFOjfuHI/JxYl3Yo9
sRX1M9XzC1AJCxbdm/lijxhhGtYyXchxTG+XOOfBLf5Kex5OjcAFAAqe3GceU2u5myrD7VQRTBA2
6r9DbX4GEHuOMKDogHaqEIOsM94FhQFWHCOZSCv07SCN037I6+qaDJTAVraAgW1oM6XlJmS/G5Ql
5HGXIlyD/hIPT+Wl2f3CvOcikBQMUWmSlrBhwsAZeFkJRidfFAA1lwQtuOSQR/k0Txx75kIDieB6
nVRtlUwOic2hapkDZYMSTQRzUyzhDI/kNAJLgdOtVlBQDAfRDk1wBBag51o/c+ZUcyBuEp9b/2F1
lQBpu27eF7Qc3nF25IGdqM3rbeG2hWPnEe7K43/X3srkyWl34Lk/V6kLKrnSR5s07Jxo2pE/6N6q
d05ZCZPW1xmj+0BQfHTjfETECIyeBFvtDqYMoeTlPvnNxWY7cFlEj3MliLRHvEq+kec8zp3R0r10
8v4GUdeNaJCmW/BQQJjuzu8b8IjCRgCVP0qNaN7oEOvaz7tWfdZ1ahZbtrK7WmOrFg27IxOUB2Jx
vSZL1RLPJ7Z0o9ihKpQXL1IQiGCbsQ7ZEWK7ZNz46JNpQSg1cEydF+2W7GFSqLLiYK4QfgrbQhZv
6xQcCwqMBqQJWeD23P21BuyHwlYz2QzfsnGmaZRvv6rL/8fBQ/9mmq8+adKvir/Hmdzzovyhv1AN
Bag9jEBkAWXRarMV1GLhtJn981lrBSZNWceyX4QeMN3XmdyNo3UNf4VE1z4uenAOAzn+2fFa4rj2
c5M8RXfWoyr1RGPvtn4oByu3UYirFKV2NRtmABLCgEWFetUXeizFsW3WoVwujM7m1b+25tVx/5Xo
i+EFR7qyi2VnBqIuw73QTx3eCMTXJKzzH//V0oyRpXYQ9uf6vBf8tsYWx3J6oYj6RGHi7p8h5LtE
QdrBwXVvLRWaT1ES/ODzIdfZgCJu3Lnvek1Jhu60MN74Cgk9by5dewL1g0EpOczDJ8fh2I7GRhw3
AlxeloNEEUgURfDhyQcXFrJlEAU7ei3Bxt0gz/dXB2T76N2nTDlLZHOt10p3t4q25YU1BXhRjTX/
VNSCmWWWAf1NRDmViAubRGhpsC9iJmzYzla0MPtg6r8SMIx4C2/i63W6HkvGT5XAl0hMrlHvNnFU
hKj1yCy3I+ILCCNcbjNh1KD9bsaq691CoB07FvY9WJzBl+CirMLoR1EiFCwTFBd7dJAYYPOpziBx
NVtYxFt4Xh2Fq1dXlQqUmwoxR2huag7r95JK4H33EuWEAim/xo1Odp4zckwG8BtKs0w+4aPIbAXc
vZdGT4Tuq/jvel1sOC3Cj1Z8kfTe36mJgPhKnsbxQhDJXfCVjUXRuLcytc1IxQ9oByRtwj+wk7Jp
45puUkgtsDyM7Bjb3smXsTnEvpGpp1iNPaMTFhSfANsf65J2099Azdu+B9FPbDlHraNhtCe5waaf
34bg9yjsvWHkRjdj8/FU/tMQpZzfcIkCXADZeWaCin5dnuiVGh911UmJ6KDnZN7RdK7QQ6MoF92E
eaHSnCbrbW2X724bCfGg3ZcnKaizjvDQ9SRACtWwNLMxc9y0J/zeb7KuIubj7f8fl5+3dBIqqcEB
p20nZ4XbzqoblpHEkMQiBmSJkzjZ71rv75GLKh7kfaNbXHzu2QpB/fH8AbXvbz6zVdsnWFZgtrCO
rmifCBR10HhrZDFObIL0z8vFo+sWsYnq2+dVNl7fia69pwzC0xRvpvH3C5PD7zAGrfEiOnocI/9u
Z+iO4L6VlDWXxUPK2v7QPb4rXbp1WDrrb1K3Zd5u2v+YRsA2lWYe+oXqYqZnKCVzvGhVWFwZwyYt
EGu/qmNG3ShAxiE5O8mxnOpzueRnV/3kwFV0vci2nARLighatmKRGMRyKGUPCyhvHi8B6cyyaqRC
fWXjjFYPp39g3Fj2x1o2Nno9AEMRlLHzhT/CzmAzzFM8b986ZxNkvBARB3FtYjNOoEBSOTI8KeAG
VPUgIqP/WapEIFVuteT0H/eZ+JxhYIDB1/7LOPQLXUAecmr5XeR4w3KGoxZTbVO11Wp9i4ciUbey
I6SvMvhLHwKTMOQlEFhuR8m1Um/dNNqwGvOoCetPfZENITw3vh9pstVflPeTIaAvS9ru67kSIwEh
UzYQzUAsdYN1jduRKufRknIhzjZYM4FOUyzvz3XZx0v6kZUjxX1ybuZHIF7svhq5qJshKyBRZPRZ
nNeNIUC/2MsDlwi4S+axxqtJRQ1Uuiw2a35YXH+pEFWuPC/c6UtVSHJ66aKtDFCtvq74lkGex+sn
FQ6Bvicja50UMvbEiPSLHkd/oDl6sNLIIz6jf01LVN1y4+m6hzQpVG3gDiKygwQ56I2ns9Neh82c
DMSU2c10bh+OiNra/EOknmp1ykWClgHNfnGCgV3YvGOqDfU2GRurBGVtIj0tcn8LUKTwP37TcGq2
t7glnfrljEmUB4wnmAaeBKZsvWO3VYxMq8GifPh7ce6T4ZGYXu0J2KTtp7/YP1hlkbnFXHYQwIZM
uQIKSB2l5XCAagDPOm+Ty5HHo+YBXPO7cKzrwOcU/LEcE9ebLvqNDZdGdLwzb+D99jVUlYtSuMxu
vB0YEz60qKhZZUIARKiMzOzc2WCLxTT2Cd0Ufy8t9Jp3fGsYYzZrOifGGjmYrl9libfGTF8M4s6a
sA4wjLUfK/yskzuoA4berswBsIxOk5aVPCSe71gm+kAgV9wIWRXnFMEpkgE1WtxC9ExrBwnVt91O
Et1yr83XbDlOUl4+NGb1yDdcduHfrr/SKpaPsfN9N/hxfXJEbUnoN0gqp/1QaVbTDhVe32Wy0mns
Ln5w4/1rUyaUVdtn4HWgFuK8O3dTgyt9MTBmMKXTBBfQj+ToXPpuNyeC9vCmwG2sFXZNqgtQRT5C
syaKH2bBHDoAlT2NJD69XlO4PlLHHCAdWJk+Kgss8+ikNuIAXwV82qelWCapSzF0UGB0BxwEjuJV
dCakSOL1Nj8mgQWTSn7mL6xocwXlLh4DkIm2WTOw1FDjM/4eGcEm3gHaoRcLCwtm2Sgh5++Ec15U
Q+hW41ZR9O1xrAp7Ys4c7B3W4SKGv2k1399Vy06aKYIkobjpL6WqE52VxOqhBbrVZdeJjDTVf5BX
Q3mxURXalTE7/506Oz65u/0xIjEHzcAKWDsMZsdLNH6+Ic20T5sLIVdnWQKoLpjiH01kQ09N0f0y
sXs1DKFewu0XR4B3xGL6Thyd3kiuruwWhc4b+OOUAKhq3e+p9d9ZGj7O9OsgvbMRHnKd3viKFudK
LzC/AYAJefZYiKdYiGsNlYkFDCNCUxLHN+I8MTLz+gsyNGdDDqAj16e1xd29QrEhE2pk+e49F/e3
KIEFOYYlLo1vXVqlSHjz19mcRrOfS1y8Xm3TEMK8vqUvboFIyEp9S+ilaXCwFh2kVg8f9sh1Sjpd
murwBV+ienmfXEPJ8tHqJn5cmduSS+1T/l0Fb1vFRxThxeOpFtB+PaBuJ7O6u2/ijyJklFIKqtUX
Q7tnyck9fcdrhmV6WuHVOphhImn9Rw7Jpq10v9tP7UftSB31/GyPRRAPZW/lsH2p5NeXxhMRvE8q
2BAXndJmhHefISwEnqep0cb6XP5a7qOXMS4cfGJqjhLv7ZuDO3U7L07t7I2XiiNmtKMa6r/my3M9
f8FqodcKrKszow+l/gSAvEJ670Kz/LJIwmDxXCDEMeb3ehcdgQLEcAjVT2ccBod3mIE2tVH28VBO
tndELgUD0GPbkJNL333Q66WDMyVn4uCSWwMsbmYz8eqSFNESOWcZWcvfGbWk6Qg4fSRFqOSOdApN
veeZJxBgOW4CKONWZ8oQF+DQH4KUJ6jHqrxBfEZb6qrN9fb+n/8h67AqD0OeQ9sykpFk15c4QNr1
AJCElOMkUiiVemycF6GSrUZgj7N0wtvrMctzywyYs1D4ONN1TbkwGLt2PpKQwgrRFi2B98wrxFEf
fHeE3XfEeohoguEokjPvLybIDB6MbQQcfiO679dsQcjjoO+mWuyqFau6poJF82J/9eDQ0mZD5bp5
gxzC9FOGb7Y0PtVtCwnRXq0WvvtU0HyRQ7+RFPfMHIKd++W1ixswsGEaoC/TaKzR2b/UIV/56CeD
fp7su3mKhtEOoAUuyhgcEJG4eqU28YNjDD9BvJXv6Y2OAUJaoH+907lNkMLBnHAcK5FuMLF2MIPL
wlhtHk+R0SCZoL2eFkEaErCLxkJNWIpOBh8dsm9QJzxC5i+eRxsBNlcpX2xu6OU3Jo7MC8fT4LaV
ZCcg2pXyyCe/JZYJ+m5Qs993wTDaElX7dskpnljsf92ImXh6pQgCnqdvMcsOzIow/lQS0jmv2h+s
721LPxx+nVJ4jD7bFzxxQBnt7nH6wx7Yo9nb2jAJyQtYCil9b6H1I6N1RqQGNqioD/OraEFASYsW
BMB7tQkulZxgAv7jQ1QvBsNU/SoaErAm4KJWo12UOSJmeBIvr/evYe2ryuQFahCkMS6rCae576BP
sppjDaQFGKb8uZoUeDYAATv+e07FFTQ2P6MInQ6mIsDExGta252wo3370MhHSSMtKpf2MOdeRFMD
pfTCZoFByE7vhDXOWSnbFsa9smWTWP16CfqokkNTbG91QHdb4RaWTugHF/ntkKCDpVtOdRulmeyM
IndoS8stIxBK73XLeIrDD8wjTgJBo82en/EucXPYkz58n8UnJagLsu6tL/G4BZNi8B/y9suiqstg
nVxl6pslqoj67xXjEbhIDdCFZDkd6rlojmxtHeyZSHoEG8F37yoCm5Mn0pg8tvF47OXkuC+waD2e
lj2bucWTaKD0WiUVcuN0uX8IF9nt+S5M94rqWwgtdwrv83ex6o9jwRHKBq5ZxNj+GhR2Z69Q2ffa
AHB0vsJlT0F+ydByVfNyLJMoWGsXQ1pCHzcv3lt/qGvO44N/VnMaTlX79mU90V+0HqjLquYO3mX1
6yCwVkLjrvtAln5J0ue6bcFzuUnS51kMhb3Z0NIWWzGcm3NA1ebRmzxQtEp6BYCg1BrlNcgQmaHx
rrS45Kd5iixmJyfESEIZRLV0S+nSc4U8VD+SyZfC/QirnKub1lbnLsLaMoYjE6oRRSB+K5nuVN+c
fuYkWOK0hvQvSyKQRzinkSUDW5V4/m9o7kYYkOahZVckZ90S72Cv9vSrgzlbncggc3iuTPIhFa/c
Bb/bHYq/Pv05chEOnzybj5K5BJX+jTZ1eLTwgJHZPAKhObKjOWW80sY+rPojd++Uk8VyPsSqbTL5
o1f5SVJB01tNxlfn4GmRy0Wd/kCTUp0oRHM8SU3TPj2ayqAV7pAV6XO4I21RblLrAPrbJIFWdZ39
VB5V0ALCOXJ8Q3LpRueC2GnjGi0bE73LpjBRc1aSx117fRMJEi+4KZ0h44qOjFqz+4KaRg/ElNp6
huolN5GxSt9m2gMQpe5NVe3LPTAUwy+VvEd7AYtTcJu+p/NMdCNEKGQK1Hd+axhRLTYApbpAg5w8
yxPkwf3CTnwnHoM62zuAGDfL81BnqEVwsfpKdLm+JinhC5TAi+A4q/tutryWDVwT3Id5jPCVReHC
5ZpUL31nCPj4mA+MjoAbFfzd5FU7vNmUGCe8EuF9yPbtwcNpewk/Mvdghs8ohSt0l6bTkZr9UaOM
sYl5/Vl5xaSDiHwUiGIkB3xGMiu2JOZCl42PiOVLIpMYdu1oFankETeRHkLVLWmJrqwLxjQu0oGV
MCfKjI3nhaA00/WRG24e1af/0j8ohSqa8pFyIp3NRWG72z8K4/0Wlwl3hGeaCtI3GRJWb1l+ZQe7
5HwJD4mAAvrewrkkPgYnD52VqQ30nKKRDJEWc1MlIB/ScR4YLCNjdyV38LOnG9ZTWB9JDc7oIZsK
OsS2RwtWqFvavid61wtHQkw5fSP6k0eDonSHuExL++jYaVIKGtc1CBgYes4egcTECquhOcNbvcF/
rsHJ4Jd0mTHb0d70T5fdN4c7pQwzO8buZVsKyRGpe4XTY0112tdiJpCzC1sPoX9FpAOqbih+2/To
12skA2F/JvL90u6ZJHtuQ9zQ3THUUO2uvZw5uPm3MQl5TrcaYmG8RfqvB67ybm+VvG8DOkr50svf
0+r84Jsrwm5JSLX1dV1+bwz/pve2M9qyyge+jUnk3e4pluUJN2DrM+JaeZny013yMeL2uynRbORO
oMRzrrTsihmLb7q80jrYJC8eIqJvDmjtpYqOcikY1uvnOHbTmy0G0yLSwmM8h1of+d6BzJAgj0Uv
UxfXgeAkW5cSQ8u8bzwae/thXtuhTgM754zpvGlyoGAcKv/IfrqoVRzh+GCXhKAxBBH/hLezkfIh
/VOiEkOeq/RmaZMSADiBriWRvxltRb4+cw3Xxz6fyy7V38DEURKBNWQeWl5SjT1r12bakhV4NvBj
GhLJIpYcxaMtj6diA66nIn2rL1h86Ldxvc1fH269E00/KPqI1TqoE14NJTKNpO1tL4FBy9ReWkrT
Yq/UEq9jFEEobflY52lYJUakU5hbS7qdBbPgnJZ0Vzl1BKsSaWFkHYmqUYwOOO1cnRDYGcNavt+Y
iIv8wrH/AgesnPqVl8gJVYTIf3liCzjJ04xycf/8bpnAg5NVGDqvSyvAN4A09krZT2+UrRsYw+Oy
PyHmguUgsgXRGMNiF9eFWwIhwj1rT5SQAyO3u6gYosdO59GmpiRexwPbjwitiGqwSST0X9JCj/gg
m/9m2Bl6bxQm3Ly2wx55r13NfsW+rqvtXxDcshAkEWCPE5aurkC/i5PUoYRRnPUNRfbEBUY7/qg2
UGMr5pSvsIqML5Gr/7QQWoGTAg565tylMpqne16gAndlUuq2G5DRBHLgRTNQ6PNQ0aucHdrVvoKB
DRTIpWKMB5r8jwBZB2Gk89esdLqzr+TEgh+WmNe6h+erCzH+CHbYL04cpcourANQfNxadUJn17xR
Ib62IY6FSGA7epoxoR93teW7dywyziYxyYMq+/oywL1XnJGhBFYLwXjedMTdreIcDbkidoNZM+0y
Ke80rJVu+SsD4cPTCWTmYBs0kg02+W6nMWzW9XX9eS4jL2UfiQPhpSU1GgwQ5Gia2YScMB4YYp6g
z0QT7QebRLhOT5ukj36Hzjrcx66yN8aQcq7sxeIjiGnPaHLPgY2iLNtlwwVLvn1dswiS3quklFin
THK9p4j3zCqZ7XdH90lm7dEbleHSz96gK7djQNGE4e7ebwXqaUl4FHupXxCnsUuMCTL4ns8KGYL5
35OmDaa6DxMYlNztrwJ+jUi1P2sPpm7IZ7/Z6DN9QyQcT7Rh0E3L5ZW9M8KZX6QsYDV+T6GXLF8z
pYcpxcIdrT3NfWLv7/9dNX9YHdamNTMncGI54m8//gWkxj6yhTC5Wv+n7WmIQeBno7d34kA75c7d
EwQvMt2pzuO9tUA9k5kvDPNF9F1QBYdGzPUxoB/LMNUj+jfJSPoat8hZKe1rC9NmMakYJMmmHmAi
aWDssSoi2Qx7S85vBjz8DnYeCb/W5GKWVLjAGS9nZ3bd0f0w3PQvSzTLLx11A8YAIW6fphl1f0/M
ZGAp6yLYs3OM+zcnVH9i6qEgq3TmYwK3WVOHboi1uzId2anTpJzcNWPd8TS1Hdt+zF57qzXMaM22
eiHVNxLQaRP/QHX0pDTYl0/JVWfKiTV2l6Gk6fzSBQzFPrGksOMNVNWARYQiW2G78Nmx7Mhy+ahJ
fYDybqWpmjDw20Pa7DW3dX2j+cRqw9CZYRRjGQY6IaxmFE8ZICFJGZvAwfHECiAtwCY5eCJAlC37
0iSrp23/gPSCNdeqplmexNPEv0fkstMiAWSrzib6DmDMG2DYgCnYL0EjvLn/CpUeuh53yFF3xdvZ
q2thphdS8uTItJdNVW2cyeYMMzqsR/DttlSe9+/Fujk/TfuFdqXhr2GVNZNpR9bXCQxgXmZ/BpVT
HAvpcHBEr0pjoUDVxDXzAdyNgQ3VG1WGsAfEORihIMxNGYX2BeHJOrE3kUFNk3kMcbHyzTa7fU5j
zXP3CoKJwD2EbbzNijtOKQALdHrjL27nadr/N5UDHdVHXBuXH2H2vFfJHQZbs5BZ+9xuT4Fh2aON
gSv9J8v+WR1FLORzojw88Rqs2F9TS/Njfte6Kf/f5LfZaAfqDbf4rH9VxDlQIAYde5ZJTBWZGvqb
l3w5138qnSXrcjUWtp1JZKLarynVtdkiLuoIWha5qK/1MCkPY3swIzJyHPba191g9zblcyw496NB
EtMHCfZ3vgXRotHXeW0n1itBApfO4+BREsh30Ox78GDno2p1X4MA65V6bVgRsHy70VoGzhsNZWlt
Jl26YB03eNW3Z0t3ElReuGn3WGHyfmhw9xuesRDBexC6QiK3WyhKVCYwhAFI4PKfseAVzm1pEijo
xm282ApbW2U5TjhDFuMr86J/Xjz1AX7D+F7H26y89LSMpN5dC6JQCzna57nmYNljMZ1kSzUWEW0H
MHPXFvF2PH7jQivgcrZFCaLc0ZgrHbz4Pdem/VkTlrLyINpWuNCOhG72tg0wSEcEP5zCFeeMKKo4
6kllcsG+o+gGvEfheFafxJFbqhIEFY/Qo5cGjUqYRcogJXh3forjMe4LKCNM1uYfllhR7pqcr3MG
II8T/daI2aOsPAgz/FXY+XnAIOs9uRRg5aJsbqIJJCQH6qaEf2RL48F76vSheVbKTzexMryAiHCx
rc8z4qvYBmINxEK/vzru9+edW5aUKRw6LAf6esKrYpEudP4GWdTbB6Mln9C1Ue0le71/Kr3Pmo8v
2qVTR69SHsKDXcky1/8LTOJkWNpjneC28tO69ks8mtErDQL82AKNw3jEwV4dWjKA+ETZKWUito/h
vgsiOGtACPd08VCgdo04WhuNJhp5z4Swv0IqkpFE0BzHH3K//0/Yl1Z+/KjCbtJY2tlVmT/ow+Zx
+do5f8eROb+gmAZlgs6yH6bnMnO4QvnrI1pjGZHSFV+aIbXgLKThxFu3tT9Yj9SuSjWjauibKUG8
o5l3nchYDxAqMUFGC/HNErBUAi0fx21ji41AlGEyV10cs0abtnIa/9V24hPmvnhjGipZW9ouI0SH
KDe5Z5/xv0qAqGfmm0jd+d/5X1gD2mRQtGSmqyIbCH/+gUT0FTz7dfaKZd2NDVk3MvACIJRJH5oJ
lEismhd1j3r7yIz9uKPOC/8qYCwoLoSDd3rDf22eg1o2HSzr2HjCs3sdkl2/dSoToXQsEzR1X8fN
XHvOUURt2+f3lZGU1W49M9+6W754QiD38CkLdEKOdeo3KI3icl9XgdhyXT/uCoNuEcH4+vDQAgHI
pqsD8cDTCJkzRGMjCqSnjLYWqYC+QRhNCJBoTnwZIpeDca/wf3HafIcx8sAOwYH0Mp3C9oiPS2Wl
KyPCmthfgo5hOlVicRWJUU4lUuG4Z3dhgW0E9mj+J4bAijmXCzxF6I9OaSy7qB7yQUZGjpq3Y8Yv
tfRMUs4AnKiynhM41e7XdrfcTE4fsPctiG8n0KIw6JHMRYOYY9ewGD5bMxgpPaL8iQ9vdGianz82
Yf7Smgy1WkWFCAMsaDFf4lmBpnZO/Ab+Jtl4dclcOzK1+ccDHYcdikPS9XyxEJYmOdOfgodHKfGE
o2o/Gw+lMLkNCnu+67iOYHfDZcyIzXMVgXUsdEkp7AgWqvTW4eLZQCIi6t6sZye86pdPzcGOHaQG
sY/QEsbkZbyVsVl95N2hnuDgQpeok05MoAUPOg9nyeTwpKwDjVqHf+x1f690ip4m314dDnAJ4lUE
9ku4JF9vhaHF6W+mB4yeYof2YkzPZWjDhbhiT5jzxM1K+zf6itIBm1LZODEs4s70hgyWFRjid+dt
l5Sj6q5bqLqOVl6GeipDKOyCe5VuV5Bu9P5mX68QTTJ80PZaU1cLV62xBw8j+4vLJA4vVicnfT9m
sEjPVJqm/Z72Y+BRYVq7ut3grp+PGRGg8xbERzfIvu6xJ0Vr9v0WbHrJ6T9S2PIVI/5/lCyFwJWj
luXBAd8EUL4D0E0xYq7+CMaf9LexYmuj9l6YvcdOFjBuLVzWpjaT9KtOTnI/AelrFP6HIfDsLd//
7ip9deuLVmwhe6hfCJ76I9BzcDdSx/mcou6hHJ3ePJfnuXIl3NmNIwhBT+r6E5VOeV5e4E5vBja+
ZgctmRKc4Ld3PBpdJoR+q6H4ViF2onGpgyBu2kejSyLTD6TNIBewlJJI4D02frELuIwJt+Mnbvrp
/WfBiTABM6bQqf41Lvls0wqW5XoKG1QtDNmf15VOSDnqDIhvcNb5vyKxssQ5Y8K01FZGABBUqxXg
z1gJ6I3vyUoDLfazyxSrFVTIKfhPkR8fjEXt55XFIBhD7jP2AnwFzvWIOhOuLVtJSkIECGvuUYM1
Dnrfv5wqswzMMZtKQNI3fs8I1ISimpTpnR/bp7byKLK9bxqhFGs9n9LFHuqrRWTBaH2YiD+/9t6B
Opp+TopdKjW3o37hX28QQkSAcqK7JnaOAObxJIV4sSum8bPOCScL+svioh0RoDQcRiwfrU63LyZ4
mYCAywUegQH4w36U8F1g6q6NFYRXn7e51k6zEDBlZP8agal2V5ZDeRENVdusTduoDzXVKWOITW5b
3L2HXlGj5cOcOUTOBXCfP075GmyEozca22iur4hJ90rVugIqUSkSFdB6GjllfrFsozqCJKM/w727
NwlwTAQ9dIIQhJM9Daq8QfrdwaboUubuJ2F0F3VhRxzBtyffrs9Qh30Gc/Pg7VDv9Qip+p0m+3+L
x+4hvC2A3e+r3US/5z+6ltnMAt7twq/qI9fMNYspVlLyGmbwfXuHjvUYEYtwyFOHIsAhm38qvK9O
ifJSojieovDVmWm3zCxJ4rqZiiFiC//lK9VR1QSZsHuQYXGUpmN8WcLxOK3KNMTZbUIrTBBEM+8h
WVu38elpb45Pb7OK5NvIagW6wRn++N/GDSg+i6PaV4uhBiTdnmQS2pvfQw4+W57LEI8FgYGCNz5u
jRrkQAFC1fUtAiSUnJ6q1zKxVV10lK5Bq4Zb4Q82ekrI2kZYzJLsLNTFglgtMLnaGltfs8QQR8Kq
ZVb9DelO9mt9JwuKfTXElXjJXYsCDFPtMEhPXb96MyC3r+3hJi/mr0K2+Zfd3ndLQNi1eDlRT9PY
5seN+Qap48m0jIOJ+xkuFhHNavufvlpJ9xe0DxHi1O73wP+tUAjkr+deGKbw2HW5RU5nT9hifRF0
I2/q6mg/M1n1z5BdqFJvu8BCoQFsizoOWNNSDEK5WTupfJhpLxt1BcRCoxNNofiVLyqS3dAgtDe3
wyo+O4gHXXL9NBeGswt6RQ68UIYszoISOUsHCr0Ry8PeHNSGNrh2yogkpABkFkBfjYlWNaqu2Keg
+BV5FPSW6Pw//V/JErhXxqvkmwHMoX9oReWVb2wGQ2buO4NXxWMJLvEHYwVUeBE1pbEIpC029ISj
Q1QP/Em310bbiTmnStWWR1wuv/itbX7bHN1aDUbI1ytleaeEnQ8heAZI5+X20iCIcvu7ohKyXoEa
7wyXy8xEFpgGbsTv/s6SvkOzWGkafevy+HbNWZcgV6fMBtUs3kzmnvXGr/IQEUJBP918WRob3TzT
PIJZ/QxK+AS3r51WVkElBiDJj3u/7ioD41IOWZ/dGhyj+FXA+KZtn1N+F+GKEYySVm8yqZTWYbvX
jLa5q6ZRhNB5pL5j2sokR5JuHN4h06MzmAI5XsR2tEzG+H7lPtDPXf5eS0sTlvVZ33Y2JNFrnh1R
LLfeREZjgWDG58wh8CNCaL3QPZ+4s/CS7K0ZPzF2VUjE1/22SV1vdob9XVp4iECZLokqELdTCTjG
nuRMQKSaFHo9zBVfqD8H38nZE3DCIxAplWlpyQXK/+hgRuWxSxLO6S4j/NObQx59lauXuWbhZl8r
ATI8zDeJmTJlWdiNuxg+mnqI/z2FLE2kmX+Tct8IlTtrjijMMqNiuGDc9Y27zFKDMKS4yCcXtzqr
nKiC9q1OKeydkHpEzPV/Ld/fCfDbcI5CTVTas7I1IM7lrUZUwO5NgjYJwSXHelfsTeeymbzvZ1RF
bi6pubng246BILe/wvLzzkadGFw4pzIBmJd5SfvG93CGzceRnKcXTJ5f0nZGK1q2Q/bz/Ehwy1GB
AsBRO74s2SExzNPW2UGmj+Z7lMVeoIg6dCXDe0jXFU8ZBU7i5+KUXNsJ0DC96h1L6ivV+cQTGtY5
WN+qWKGoKMkQPprL8lc/tz0t6ucXfTB7ofXIlip4GcpbaaDmbHLBEO8D0WuywUVRMtJKQYlhjWNl
qL+S2TNxv0nW3p3otgzsPcUDCIbwrkUlMuz6BQsFp7ewaT7zlmZZdctaP6wTaAqj09gvcF2K2nNN
MO7WBQh4lDUjY36zXbqI9ajXWutIdFMj3xsBFbS9pGPq2rOQoomf1FhV6CyyYBHpF/GJtrYuulMz
OnAmgPyDNU5R2iWFFjHeo4biJkUqwci5hkc8UXOxfLayAljl+VJ46d9eq/msXTdHO5wHiK+ffKbr
5mWS+PO35MEkQCq3G+7UpFUUQRWmLhEPsFda43mAcOAMrhmv0C34DNSK0saUlg4JZPH/gv3zTBYn
99FR1p1iaBaXb1sAGgWbrwsu+EuDQkLmwCxzQ484IWjEa0FUD4f2slhDofCTBbH962CCzd8GSail
EuiXEKK9q2OeXOf3aJpQ9u6Q808VhH6/N8ZPkHb7RfcmcmrqmCoIT+CbTGUaB2+BgxoZNRVa8xc0
xqBNC9PMLSJufOZX+Z9FXQb5uRwkwTyQtkj2RDl4mtLDODSd1jT470is7ZlM45lhK8fUxHacAcR3
R+VTn7Aab1KYEn/JgHJSp2NHEnGNKpLTQ6GtGf9fSsycGI1wQMRLSI+xBFwUWdOXcQy9zCvMy/Yv
P+SH7im+V5lx7pkVU1WmgW7AL45m6uERlwmsLZTMHSI71/X0WH6n+DHb6xTN0kauuFvAFXiTX6VJ
jkjO/gLLVVSS4oPzdrvrHNqXIxpsVu5/ANW0eQOiH7AmSThX9JSa1+3Yx15msDIG0iEj6IXoz3eL
PG2bM/rUEhUWliXaXsMSr2Eo5dPd/gkXiefLxIFgQNf+lTF9WxdsYUE9Xd5yhWckRCL1gy1VSdr+
sB7niQbHKLkSJJKUVGR614Dy6+aQUjHQnw+78d5rjzc1XFcU10lM4KRywuW4c99Bbph11yPg6A1z
coZFUb4U1Hrc6OfBNHrseTNrzBjml+TYELoBVB6qDwtK+7WghWO5Qxozxp14AcqE+c0BTlL5lfLg
yzl1E87cMxAj6YwsCv/4eOzeMpnW+HMAMAvtCkb4y0j6rRB11D++Hq8hn0of259ar6gG/xJmF4nQ
7nR4yjjfqczH2rMYe4oOqDVl31wMNpACDY2GtkeY0mtv/AESQdwnJcWrMygd+4ahXepj/2UhgnpK
EyJ+PmM3ahMsPJiZGv4g/wdE99V58dUYFBKyaU5N0al5bpeQWEk/KPoodW1vq9y3lvXrLGNDVQnk
M5ACWG+lwRT9hRQ927zmWuv430zia9FXlmPTIh/NLvosCEHUiX9yvsZi+/ororw9c/Z9shIlurZp
4TqFJ2x06Ga30kWX20DsSpwIbZ3FjM2HirO4w8l+SdrLIsz7znkA83EvnngS7yBsBzHFeILFQFCK
9FLRHP32V/vvRstSul+xUl0SMT/EVBIzrI6HCwbx3x1c1ww9pXFCIsi9/pi7N/HU3QAQe4lDx3vT
5ohdHym3wp3O3gXPZIyzr80bh+Mx9Y7ClTPKke/Jv/108HxluNXrIGthYD2JlCiH67Y83Pg8WoKm
q1mKTW6zQSmG0Q6+zxjCnF/7VwYrkzAdmFILv61OnJzVZt1MBVh5FfxUYY/s9zi/bs3ufarjrj2f
mnqsQtqcdTpmle4FmP7UdMUI4CATup1NT2Bs6N0iVPGz/tnL2iAwmLV1yGgxjAZSsa3rjOCBGhqB
QwVNG2kn5MoGqTgddHHcfFGN4Uis72OVehrqXBflxMUkvjaRkDuyCerZjO9liouJNh/NgCCd5ts/
/1yb9L46FiyEoSeWia2ExGqSeJs3yhYgEo32Piin2SM8N2RwgFqaWqsPBYM1l+lITZPdr0Ooo/WF
bfrk3YesKRbUal5rqpWrj8PSibU9DbQ+ccP0zdAYtx0ukrivMs69yqLqa8a0sB5LofO7jeddPP4G
W9llv265GKK/gTzybIS/5tfVEjRJjRtd+Qsrb094+314/9+x5h3gVd12JZ807EbYrLUqcn9UyDZW
y6JHV8sVJBryoYwQ46JEijSxyZkAIN8VjLXDTC8A0OHYbdbGDMAvwjYPxV1Es0ybYr4xciEa4NkK
N20xKJiK07O6KBvTXEOahasCUotYH6G3Sr+1O5qYSpwC1hD7nS0RzOPAAwnp28uHZAaTMO+cIxbN
976G4q4fw2gC+czWG8Fgs8TSt2UIWg6H8+QXOTxuM1axUXbmDsErIYPz8lGiRKby1MW2LJKOTpbO
y9Mq3b61ngs99iDmCR2B7YvJGeKoZSNHdNgWzhyT1bf1oCN5vKFz4SbtaFGVP99N2o2LVlCwTZwZ
IEDNJ34a5KKaS3r2Mtcnj49vqabe11KZ8zj/Qe4AlK1yvOhKKcNFU8Xx3Y8cEqdF41X+qGIhxpPx
t/bOg+L/X7SncL/V8+KyW+7MV2Ii7b0qeFVtN91GbdEGpoapuIvvmNOXzKjt48D+KmcvA8JmQccJ
B3fgIftoGHALzMiNvCdfXijdseJ8GelZEru0Oj2VaIflyCQSGTANcc7PTCZdw0bX1H2kI8vUG/qr
3sQ4X6Hlh0ePwxg8NsQzvg7SkVD2o3fwoQVOg3p4jQe1Ia+47uuz8sHciFI5GP4dLUEgcobb9Idr
3DL+otgij2KSH5BgQGvuvfFyOMjvRJH2ePZmgg+IrT0/7f6BrnZU0iHFlIxJd25JYkLZHLl1gTgr
LE5HxMh0Q5vKgbVCStrRERw4XX8GwvHFhOe2SoNiz4QhbbqDNWucBxj4v3mj6qEF7fgmyaESmL0f
5mz5j1id+Zfpvgb9P/PR2WzJlQ78lX74iZY5Yn0AnzOTZd4BLcwDoqCwbPkJPWPlg43r6Q40fXHK
gShGevle0iUha+wqIe6bfZWMkIMJPw/LVpx4UlV8wMmxGuSMgW5K3Uub523/xHKjav++IRi+LMyy
rjQFoBN1In0MFOI9HEfM1Q6oFUTVRtT81CIrr03zhCC6CZs8xZELUf0dOrAziKzVQEe0dvaed6nP
L9OiW5vueaOkF6eJnxJJoLgnX4D5ACva7sVTudN3nN7lrOMIMPMSjFw23eQeY8JmW8bnBFgJkYb4
tGWdQx6xK7mKO2stRMOBO96HTjkvkyMHUb9RyuRfI5tfXk1J9lsP4Rs5YUOgYdp+MdBmvUWb9oek
FldrolZcq791UHRLoWtDwBBnyETSV7t/USTguT7KrZtY0zsoMbM370p/clCH5u6pek50W96bxcu/
WLg7UpIaZ/R1lX3MWJW32BVEX3f4+wyfgxIywXVPHWucxROq+YQ/flat3tVzuxZN3UfXyGceDcmL
NfPHEDXcZ4IRZLXCRLZvyYmwLv9MjziqxVdavsjJEb4MYOlWIk92b1H+NKJwu8ucA2shOrDTlrjS
MysvJ6TNU6sEk5rF2bOKVRh5uh9cUemWva8tJJ1InL+hZZnDv0iKYY0HOz8imnv2Eg9s4DYf6yCV
WjIhR4ZQuvBO57jUpZ3fBgop1aUyMedb/PsZ4k55v3K3LudMeZpRfpHBfeuM3BIcW0rcqLom0zgq
N4TIqAPB+gW+Ah+75uMZnWujl9SXraLuOIjZvUL4beaAmWZrxSpx4PxcbN336N1+9X6MlkBgZITR
unLOPoUL90h+FtZjIrnILNI12PlegUj1jPObtBCS6gt5VvRiwq+QyPBDxdRPEyNtLGkThsEuIFgj
CnG33xrwGMfMbcQWYhdnUyTLJmbSPBWPQOU8oI4Gsz2cFb5lReIoiqoPU4I0DmTckp7wf3ok/BrH
iPjvUFUb1TEgXkJv7su7sdL51g8Sv8lzvmqE20WKUTXkyBIOZ0KoXeS4U0QlpV2UbI6t3pIKSv2U
0dQc5s+3N7Z6oL7WECZaX+YrwS159tIY6cf+AKeIlbrYtLL8dgmyk/RVT+y6uZGy0+GRmSzWXam3
OJcuDiRAVLnRy3ZixaMVsiN+nEVyrNA8yJ1HKRHK8Edi7/14O6JIh0dDRr7nLUCYcFWEA7kk57CB
sM1moFnzQ3VYFHhwuGBkHUCTsnwD4ylK4/D4LonBO2lKcHRejTgxLVVn6KvbYby16pUyyc8DeVtR
ghZb4AK9v3RU2FqRDU7xDxJxVusetbxktZ/9JTuABJSu/Isie0ATlOOJIWACTUh8x65vIKrFa0ZS
eBuCOqfOGBq2S36XZ6D4F1KO6sXQqw6hV0gj1+KONYIkRBJQpoR30hX3Hi0kC2z8Uouh3V8REXf0
ffY+Xo8Pg75+lRhe8d6brtBBoSqj0G8NS30W1+VuzswATW+k+fOE3dMLapMYK7SGfBwj5rE+x97I
UDou47hL2HOMA7KNBD14BdkWNU3x3LuYW6DVNp67eo7FRI8Rd+7taR+w0/UwajIvDE2dw+qvxI4V
OMCChjlmxSLKCNvIoH0hjjLm4ZwYlXWcqHPfiW681Qp9FyoYCHaBGZTlWETMuzDESBkgDW6aEjet
orY3RVUuwB64NQ9vXeuJU3UW4e+LImkG3WyzBz5xdhi1O9CvtzuDbscyTk77GoQOvcoCkEGpD2m1
itmfhQ0w4v4YBk25fU6zFAlplJ/Ny0eBYc5BkAo55wIm+iuOIlokCWyTqMV9LS0DeVfjA02Xv7YS
0+0Nr07AUp71MWs0StvR5PaIaj2unc13CgBBlcN6SGQZfJmpBx7vL0shmxF+OcgrDt7/jnp6GSro
GRzQJHU6xs7RZLMwEZ+e/zTZeB5HKr1EUsxvIMmZvOgUAP6yH5ofc9nPEA4O4tV3Ns5Wq9KygGiI
gPbSs3G/U8Me510xqbBfAYG3APaOIT/H0S5gXDr/XDVb5EfD/NKh74G/pxcHv7RQyeuasLJQjhQb
bx0Quo/huKMHo3wSA7b6pgqv4qnoAh8bKhb0chCPamx09sKbnNWkp6ekkzZ7lz1tmfPm00IdGufG
189g1EkJHN1QItT/EuFSyQ2xOAikmC1h/wttuJ5sKIvIC0wOU22DzWaklFKBMP80B7/AHwIYe5BM
fnS/nh31IveNxl1T9UOk3bFuyQCWflrNDpB5Y40MmfpXQNE7WTMyUhXZhVE5qqmbxvTxZ6BM7Hr1
FvzpFmOv7vwXTTANKI1nGYavFAQ/Szsuvj9WzKAKPZgrMMA+FhBwfrYLpnbQ8gpWiT9yPtU9fHKb
pShoK8EcGZNeaWMyVdaKo9UbJ6EobhdvwMXHvqceGWkipqH/75qrKKfJtrsFGhi0sFnODz7WmtSw
jH+mHd5VvOm0Z6gcnmu3od48SnKwEimfssYrzw1XBmv6101Un4/aJnRhpsBX7FE8iag7qVAvtWuk
nVkm3IozF17aYEi3pY3saMZGmM83XK26O3eravMYoVI1hQgBcKxapIqT6KzJ1IjzXHKjTZnvgBO+
s9/FEX/8j6YK/dadG+dz/GNRmbCcpObM09S85WKnXWujWmsLI4nW4/ER2lCtrmJZZALwaYXF3Tzd
QOLhiSrwHCf5LadSpTiqzAP5Np9/CaulT+BwakqEwI3nXoUg7zDu87bvuTTyhIb1i1YvYnDkM1Gr
28Ja8S4ZlYMO+pRj1XEOJyyGNNxVfZEVj+y5/zRQDCsjS/A6FGhHpgqkrudSqRoq5jRzhhpgaOZr
umgMWDvG0mFbY8FdqucACjZh407GcrbHsLYGyAIOmD4LUoqD9GPsUfMKRxA1Zo+7jXhfPGLFvOIY
ZhPRAza5PSMcTqcyWj1A666B8PmsdARIIhSCnp8FIRXJJEtWhn1EpoDMDfZUtBRX0DF1NI7UoTNm
4Eh2Pb7qnFnQe2nYzevGEI+O06BnIpvuj89zSgSR75UI3Jx0QzHsI2S/6Rql0zPCJYQrEMdiJamb
QLUyMTBLr4ssKIBsGAVuIQiCSNvmRjKm7RhDO2ZA85XW+BgA8tI5Tgv2XlObg6iAMAhzdcBcrhQn
P5WqY54HTjA3BQRxTGzIZIH4NlswXaafOnUb9MEtv/8Rzv7X0Jr03587i8wi8gd7WkhAcVb45jQ0
slpmlJ93A7a8bGe4y/kQI6X8BItX72nf36AK3++rf70PVVyOwXDZ4NpmW5UpkaSV3ahBopYmD0fv
qaM1wF2qHdM2vE+aIK21ej68jNySbs2W/jlnTKjxwomjI/CwqtwEjYqHMYVWuN4BUOmAEqDkyhhU
UMU0pXfEm8W/iumyeJzQzIng5F+4XJYDxmvF452VcA3/zOSj0ber2g1VtG3/H1gsdSBkL9u39Kal
2EQ8R7qXuGowVMS0fPn4uFjekn9QwtBgZd4wPA2GPIERx4aQY4KXl5nrI+oF9st2hsw3FNsej71i
qDHcJikfuyME4lSiB+1AabD/YLy1vyFksbE3tjWBuOHKliavO5ZRGOI3IwVJlHRPTO1cCcpFQm7L
PUMxcB7u4IwxmDhmC52tm4hGKsB7lXFiM9sT6M8bCwnHl2EUiNaEdRxRUbbvXnFajaPkuAEl4Nuz
0K/iMnVzea5qA944Fy17DSkjdRvTYEsd8waeqI+DOW2aJmm9YrhGy36DnI6UkYTK5BDU5plfHiB7
XkGKn/NoEtg47LSwV1L5WCy2tJ/88pi8mmnYGS6QDKEzOHIuAWZsYG14AXYcVCmR+PBB48VH+t8K
66Mzbhb5Zr0LNfjFDWdt/artImXKYzXIN23kGw5WcQCXYQITf3co0DlX60ymcC+Wqf0eZCnqAWjh
ng9h9z+XFaaGmwbFrN2++MkxF0Euf5hLQv5I9T9yTn2ttzkhs97uZn9cOjFIjRwSiizbWLNYk9eE
ocOLz+xXFkAo1Yq8h7OwDC82L02/tNE6pqS5FM3u9dMv7HeLyui2542KDWy2RurOYjRJLNmdIXDu
mZQw27oD4nvk+OtMhe/yHTXwsJaCb4UTlqei7be8hzC5SRRib4aZe1q41vnlIQ1eenX9E0iLRSrT
5zQJEaI0/qK/3w5zm+TRSFh0x467tdkl5nWJeo1sFbnBFfeVUJ3Hz9tImuEvYJPOxVkIHUynh21g
l6YlR41yf7Vuwsr2mh9TdZnTf28DeFVfUmjN38J0j/qOT3FWNXKcOn6Tbww9Bqu+lHy8GrTzDAo7
oIx66sytFhiJ/qAuo7oxO4VI2XjPArmB6pl7zGpWjfyvfy61oE2/QRuaA+r0eG0l3X/tbv5IWCAA
kQR20pe+oOcKv4b0FpLk/yIgUbSKQoVBZC6YSbF1rxX764ctX9P3M+UifJB1bm8ORDNl4Ah8511i
R5OZl8MrXeg6wz/pEtVcEi7n4tjn/rvDoOE4nizfGkd5ZVMUi5U+U1KLM9vMcV3XQvUmTMYAPniq
3ilMHzDFND+YHK/XQrmgMM+KNx9lCZgS3s6A6w6atX+oomI4gG/vrjrpqDu62IeBt1lmOzAnRrA/
fj9pEk1JyzAQ6JKFO3nhU8GI4vWFJfTNCu11u2PPrYH1+rq2inlNrFI48jTTy9bGCFol5uFG1cSk
nIsoWR6xRlcIEswMuJM18TpozVgY8Nh94kOiKtmo77ek4OeiqqbRyih/dEU3xc+ZJIGPqn0yiFAR
XHuK+P1KyOCIPZEp3V6jEZIpebNhv7h7zeQ/4NDXdmBmezr2DjgqH1zwoSexPGsWTDReFTEZ+VH6
9gq8Qjz80sevUqaCFWshzzDnENhOhJq3aQLsKIHZyD1C/rIxYD0FoIuU9hwYKcm9nncTkgfa9hiI
//vMmoCbB4Mn9HcOW3ey6vqNBpRz5w+FMlTKOIe4yV6hVKU7iZmc8/6AmXRTYD9OE2qts6E0k8q1
rWlGI6V3OR3sNvSkvccp6thmYH+3gnsMcDgmc/+yFCXc48C1hW+Q0dEV3hjjQ7F/G5D4kA9Hb4aK
T7bTJESIljl+FKPE9wwvaWGvD7zvSvTUsCHM7v8G82NL3B3o0hcmsyBoNtigt91v+1r5fPA88vZX
CiEDYPy8nVC7PJHkNU0c7vtl6cd+lqnAPXFt3+5JRQRBOl62MY76b4MLCh/GJdKb6THsjU6X2D4l
rlyLqqS8i8MpgSxAUNPPwpfb1YkhtRgKhucVwoNWTExudtNt+7anLYhxxaY1gLIWlITdYTjOHrHW
mNSTVDMkXTDgUUQeYfSY8T6GP7UhoPsrce6M6AUfpDaUWg+gJSkAPPm+jlFsa92xemGCXG12UcTb
B4rCVBZEoUWMsaIgWjvB5M2E0ggmrJpBBob8bcyv3ZwjE0S9qYk4BJYEqjlw7nbsD1X5Rb6sdbx9
irsD8bkua0Z+5DowOMgVAr7QYonUTfSaIM5TH0NqIdNFC/cJ9MyL3odul+E56eG7eN1urgQp45gK
/0v52JahQEXo5fjdB5MN1F+cELs/ZfbK4RlUiy5mBnezC9qhag1bLzzRCLmjIUWAV2ZoRpnz1JI+
G2LuUgljEXNOEuoPikV5orzqBdTwkHvvNshBOqYIZ3GhCb43G9TLhqPVruARK+vlRZfNNSX5kHZs
dCWrDp5gczLouOPsYf3qkhaSIroxsWXSSdfAFGx+LGX81iiIWgrMDeQNlfan9rQnHsU0yX1Lw3RX
1gXYIazWkpeesIphWezNFPQ2kuevU819BxiBfltjZa51g0fGCpy0FO6gstPyKz1/KNbNJH9VE0vp
HhI9SHRYYgtrs2gR5+6rec2Iq50JnX/zfyIXafX6KVT1683+CDPoy20guO9GJWjl0a7wT3GQ2iS4
Ia6gVwMxSNkOkIJE1tniMfTXPpmSd2KFLpNQ9ZA/qNd5o397Mw102r0JwMkNJGir/B4uCbtsyDR+
QBxY5CIHwn9vlQfWw9yyhxobXt4F3K1RFvyet0+X5FQxzYEfdMiwGjc6RTfuj+D/l13yeySgQdtK
Kq6+Z+D+4BSy5XDK+JI+O2sxTv9akbjJX8RQCAEMO1lxGIlsCeYXOYvZOrexACpPbA5SDw7oRs26
Hq5U5xbHJqdqcVicnez6grZewxVZyEj8kp7KudEVQ+FUxX4fZ6W2b2XWIXCCEHWUvPFITd7gIcxS
hsrG/1ghGuauzhL87eMeBEayKZVEPAxVBZjHHYT2CVZn/JvnEN6d1GmDq+Qp5CpY0PM1YFyhvFZ9
uNCLH/hDCrZWZ/QQwCeRG5pU/qf8hmyn6A5LSzGQP7Gmh4bsLq2z/UMpnjpvTx2lcykUs3xYrRZU
W4ABVPlRvRoAf8ew7x2RrVBgfMdlWwoZ7Sc32YicmfNIZ1UqqDKiVW49R6x+5U1rx0Ksh/y28IhV
Mkp/mCKXTCYAIY4lK1WOGJhoVM/IyqC/9RqR7VG4+cCUS2EJGx9CVRZfxVaJqgntFWAb8MXXr2hD
29siIgvyLp7k1anIPlSqiLEj8IRsRg13rbuASCi9yF5E1204y0gx2XSdTx/t5SQ5u4QFhFxtFJBM
w8i/bM/GPbat3rMTE/Qk7a7F3Om6qRTKqfASVWTh5DtOg4/g5cCbS8YfbLe6iLUMXC80dLJVpCKO
bxxZIYUSIwpCQjUAZk6edB5bF2W2DE8UiJilZStNC1WzbqsuLb1cLzoLeMzmMv6XAqLpjEcqbxH7
UC5tLODpXtIwTvrrr7Jgc2s+rj2D4y4u2n8kff4QnP18oeiy59U/OXIV2VF+07xDP6xqoYP4lkhe
SXjl9jLcL52FHQ+V2cqo7muaMvbBbrKOXqP04PcsXdm8Jt7UD8ekG55yDt/kM7YQdIqgxaOWKVxY
n4WwSjGhAacb6gLYr2wP5y7Wv1Ss0OLTcAMT0owi6eP++SAdVNMke94CvGuXxrFJkXs4ZI3U/u5u
FM1KBnHznmkRIdPHjhtAHL/d2Ym0mpuear1eRMBA9P+NEP//f+bVciYfAA2Tw538zfMeBmkvtZpA
Zs2oQKVa8+unNPHWfWFmOSjLpRUdrVk5Wn+EtotBzpr0LLIEb+exljeTQfDAP6GhZVHB39WMshrB
M/5ZD2NB4oFSCLPnlUZvPXJqBKDNzajKTe1h1csqxCudELsFwArkfiatIWVYuQe6HvLyIOjNsyU0
ERgEdYh2MD2aaszxO72nHTCJKvGeA0Vk1RUVcYPhJgGiG93mqwm9fY2x/K3QAl/t0qAJnbwPAF5l
88Vxu7wf28HEa9E2lMc11aVIYat8627/N8iv6JsWvF2WFXCdm6+bGPS/7/CKNYBIJgbsbLSmaexN
tgklT+ib0bZfpnmKtEacNHBq3X+j8wGy8E+mMW1QLElm5HO49IfanQd/mCcMOTmPCBGvvlyhSTco
Nh13UApbJ7U+KNvUPaJSQWiIyLdxoYyIUf4Z1WF5Wtbsmhw1st4pcYnKqFe9f+UV7vlRWufdVlqz
bHHprKA+bdzcbMZ1xeTHR6pD8ubHydc7xITRoaXJ250XKmQFyhvKWQoBTJKrsFnH3zDAYfBOF8i7
Iw4WJvZEvaO35LVEjg6AMfxg6F1tR/NjnKc6vo7oXauqv1ze1Q9xtqxGPndfQtxme7PO+M0FRH3X
e9vyBufnaf/1/LIZ7ZcAg+UfR+UD9h9lWTJh47I3m4lgcDe0EjoPdCc/5TgEGHh9BfPoct4Im+d9
SA84iEE3IrpYFTEOw2WOdmkuzGdW3gtTQQLUpiWQa+Deg7xCIjlk8pAnqoZnZYX2YDtpvlt8M48K
bWo/qOC0V+b7nmD0hQroldG7n1NexgOGF09JVsDXVaPRcB/GjmVnDC7M1bRXi/rAIA0qAUAIZmJk
1FpBvjWHwLDLsZZ31pV3NozMxnLmhDqLgXTvk6dTSpTjCmN7cdBxwJuqvx5+5DLue29DYF8I4NZl
GgYFS14jstv+2bfY28vqiOrgM1GUQdNCmgsLh9p10NxvO1x5O1dPxQAkatFfhxKYuL66HApE0soy
w2YatlCIGBeiFXSX7Z9ZpMT0c3kv+pUESkEsVNt4YNjWrdq3mHQdmLDFCsIfiasAMNtsd2uC0Qir
GUMwvF+6Y4PFl+yLkZWcdRJj2zhiwHEXOQDqdVAWkaTYdTyVthyulCdo8Z7Tqvg4/SeeImKeotnp
WHkMA3ztHX0d2WmBxvoYvao7W8zmrLjZZqsTibx6yZEpUpX8dVJiyaRcZBwSqKpwkO1esHES+4i4
efdbPMS8vqMso50PN48LiJRKufnApZ9ZaGjzGI3g5FTqQpTdguQ2n5GUwvAUfTGFrredLSr/WJs0
fQFSBegvuRKWxKXYD7BjtOuLBlfzR15SNrVh4Q3KVjN8sVfICbXgoK/8AeTOwQzKFley10/XHGS/
YyZkmYiZ6nwyFlusA48iztKRaXdPgdcUg4aeA/5SRS9tUZqAr7O5krs6liq0hiI+hYRkJOk525yc
RBW+QjkAQwoFXE4iu6Dlh2WwwAbqLQI3QA4U1FLF1+hvxtGdOQIC47K6JJs1B7PfN/ilM1T0UtLX
cJbSWBSiPExypVyai7MoXO5qTSYsxAlANGeRwNwgTJfWc0ioR9EaAJsr19QuZygXY6r7hdAbjM2b
M0QHgjApKC9uTLS6sWQqHmBRRnxzJkRQx7Jl7KK21xaMlP83KYt28ZK//muqnrI/PP2t3UCT5B8T
L5DGjVQ4TblqmdnSZ3MH4BaAn6YetxNEFAkz3Sp0P7HdGOejuQgGGZtFcGWE5Qzn/c34YFhI09+n
LMi93tGityTxHVSHP/lqoVbfYy2rXiZzO5/Ity15HT1pwAmzPElvypMlwRJ1Ol36CNw3n4BJAv4i
/EuWv5ti1hJ4CJb/ozb30XVwVLBAPrTpMjTfJvUqi3JQJS63HsPRhqJ0lnYIJ1Mv1o6RCJJPjWNU
Gw5rGW6YeKRKYu/DWACw+UOw6wJfcKom4e7/nQQouKiF7m+6mHAckAotQn1FjJ7OxbpsshkonAU+
pMVW+xA3iBOtw9I5k9Xzo/sEP9maOG9EpQvqyCAKCFpjLoH9ioT0EcOuTAF3HttHF6RzSm3cdHLw
vy1Q0RbS04ZOqlNuKVidAlWsbK1fTV3nrVkLeewstPo8WDb/Wot/Ygoic1p1eMKUnv9qHuCsThJr
/YIWC0x2yA5/zC2NQcgNbJVwOdYxnpM9oJRRzjcbilxPtBsggcEfufoJr0kDM5P6rQkUalhWGrEW
7T1CNuLr+gkn6oFwDWLdktmmR5zJXZDxlqybzBQZXEx/333H76noIuMci2C5fdxJCODDSiRRrv+Q
RGyZ8vIqeT98bDfKwj6tWoXJS9+eCj13079p/xlmRQTcTBhIDcZEo+y9Qt9Wji5VKkFQUl2SPsGM
+PiSswH4HXFfQ7uR5AI1WLDGHfaOBLU2ncDdC4AapL1ACes/iO98l9EApxSFMv/Tg+yzREcBI831
ioQTt9OfSc7VDmKbe6dci2TxXlYWK3D0GTPKwcBKGzGglmFK0AV/cPmMDoBp6vh+EMf+6EpXg+xb
jVt3PKe/2NXlXe1Rbz7a3BeuCW8HBLfGrrzcPZ5liMku20pNmn9uVQa9/GgSKj5lbdK1ki4kNNEL
WV/ZU0szRvERkuRi294yvHUKilr24H3DpflXr/TNHje+5ODIcpIqDV2r3GXdmCgT5v3E60Wrjoxk
bEChae7rYDHFbqjQWfX2YtrUUUFiHy/RtBWY6KLU9G9H0+wjG0q3JwSCoIOkzE/LzNO+hIXP8bYS
faatuHUWftaDb5doyhj++vevFaV/hZh1HFKamvLL4MMMEB6TT0VMsn2EHg6tPYc+hTJTRsgXBfBX
Ol4pq6hnrpl2mzFUQ1aEUHWlRmM6hJjRALoaJ38AafLwJJRIdBxXcIm8wu4hFID2eaGPQ/PMlzxO
WFPtfACW1Ow7rnc+qUDM6sA61h/KfhzuRz2PmdurGe+IbgG/za1ISha7kPKFRAWRy9sEdwI4YA0C
GueUicUWnN6LV/V8RpeAqYC3igbhIcq/OM74Y+Hu8EyKSdGkgz2Sflxq9zHqXsm5uivMXBb48Rpv
Nl2koC9PJRlKLH0r8QU+C+lHkYv3uNv2okJyCVZzd3TyFGToWaXZ2pdbmlrNnefEsXUt1Ub/2JUl
OFTqN7NMo2EcVDo/JVE6+rWOBk5Y4N7gda2iw4aew8erq6mOeeRzHvMf1j1tIaKUQuvtktv42nsb
GK452tOndpDzxFlNrRJNZG6p61sr8HMzijfli1qrlI2s57aQbl+ollhRyi7b1vRree76BXv4Mgqk
ZAjKYbVId3YhMTu0lo9QoKO4NFJlemqKOdXFwzEspAvXeb+wo6SNkkKAHOBulKoUyBOxYSO0CLq3
8lkoOQWRdD9xp9q/LkcPE9ey51HNAC7yv1iGQvHVjV56krpSpQVpPGXMRPkW/FWWA5eotARp3XdW
WO1v4qlT31tnCuw7HM1V2+soZmP7gCNJPlkwOrGzWvw3jsYau6OSw5xsn2rPq7jMPuzTG2S4nlYv
fSWEKSlsVyaJYHSmcafxuu6u6AUlv5ZyAl8qhNjkFuadszoAdf78jJpuW4nRUNUDCVFulzvL2m2F
B/FMnlEOKyV767I8OctSoSQj18fFOqBKjYg26LYXX/kH9LX426eBjw4Cop78UyAU3l3CxEW3dkYp
rJSzQmiPmrjoyt4pJu1wH6eXVI1+bWx+/xCSAQqGbkLXo7wGx5uW84FJ+BFDR11XdXDu8+KK4+WD
bb0L0/kdpKCV0al+644UGLRt+2Etv9R8HIu37VcfM01lRmhO6s/kdsmQA96lpqfZp1wqKPL9qTyH
TMbUohIioDYTeJpkI3loSGoIUZjW6r1L4UWWw/2JHjDKk70FFH6iQc4RuG79dRh3T1mQM/gKVzcc
RhBTpIMbQJlTCDjczPoId0JOuTPy4fJhF6L/DBnL8PFTlzohi1eVqdNimZdnzmgRH3Z6gaKz6jxF
7ApUrr9Yq5BFwCqtNB+cRX92oXLgyQzt5smksYOtpvSZ7S08mjO1+8vywQhM8Y63JOn6K7Kn2PkA
4BXBuhYqMnLwIjrHa/Myz+jUMhdjOmpJIYa0A1ajLU7JsPAPFtuTOuX+sg3Gu0QSK+OLrc5jqIrl
8LOyQ8TCJkDZuy7zVJ+lCsM+kLiYSy1pfHnM2f1lGj6lV5honU2n6ilZeJNCQ4p4TjXSrBgY18kI
lI2pUYIN18nJ2G0PM1NgRmjLj6prjgRAHxX/ZNkOgxZXHhmeWUZm9O+1DXvQqixsFbSkv1fug/wW
RFyAdNWMr/txOrzJIMDwaXl+4W9/ZqXdLtVKg7dqkrgVLjVELVDKoyLk2f5HQ6MzsjyUpUU4cdJ8
6FI0Gc8WLf6pwHxGLcdF5Jzcjt7Ew5nG2WQA1WI1l43Xx5yj8JHnK7TWBsn7wu8Vmia6bmSGazPE
g7kFdX5VaTtAVJG+9uiUg6ZDFprK2ZDlwHhJrG3YtLDjGWhsaJhON+t+Mqn+Lb0ng1vPeW86dm5a
YeuUl3DEitqu55oil3k8ZUdp9kJqoP+uAzpZ0IkBrJqc21erz6YgOIS/UbIwT1x1ANxYLyYs1GHT
u9GN6LTLpcJyAo5uAUL1ukVvwrvoqD8VQkg0aun/d1/SNo2lBJtEdmZ4bRpcmsIUbFlfmWCTTfnD
S5TWXlO3WzYTL8fAPgUZ3JbdJbsWH3dxGDa/mEYIC0ZyJIWKQHWAPuvXz/LprRTNCxC0YQiaU95O
alqF212v/ZpCN2Ysh/6OczmOoQyC3Ct69TzyBKYUKwBTHvL3P/CiwyMfuuiVjrLZWCG9rbhV6u2t
r4nyOZxC6DF/nvX4/iZWYTblcRSCtZwrigkfY5iXm8L9kKBq76ecp6pxIEwlN0cXAijyWPDxH3Es
w0fU2UmqGpUGswaH6gyEuVfbZ+wn2l+IOXcaheJZay41dOorOXBDelHuS5jwlbSiIRl/QGpZUuqM
YDfwMQ0zUOPlRKKb40o/q0W9gJk965DQvRwHltqtmtSvxfF4iFydU99WIRPoJBrOmcYWRs2r7hk7
U4ESBXsR9L6U1kajh5/r0F/iZKrG7DPcmgsi5aI6QpIOm74f36c7L+3TJB6rvv6QakM31e4A3Ue7
zK6i2UiCiQ4vR94BJqFE1eqbYbzN2d/Y9LIvJ96mqWZqpJQlV6Eja+Pkqz/O2icyHB6a7S+JS/AR
VSeKfi+zCRJD9DX7Ot33Y9xgeekykA1Gg4rUm1CptQX72ZmKKfnUlEC8V0hzsZ9LdnNZ54WQD57y
GIXyiYloO0HRBWa8ewOkeR+aAYx0NvJMyYzF5DR9SZ9P3wOwK3+uR/sr8NWelTeNsbLA5c1tM+Lm
DaS7AJthW7ogGTjtwVYZe17JXLbHI3WigUXKA+BVMNPXL+7dWLeF3q8lzZgR8GCwcUt8kZAEfCx3
24oNF3ROlFQWvL6jaTeERrmvcR0eyuOA7WQy04/GW7huflIXS1JimOFJA4opeRrWZQZBGv+ep4sO
oP7k014LWnKnFPqls7niNLia3pwv+o/Lcr5IlPoCbTon+JEHxEfAcQs1zr7FglpRyxvhTcviTag/
nFNJxDAqL+i4sUsl6IvsPIoHBRJZ6ryDxX+FvOzA+WznApTFsdrYsELD3u33HIVXUxEQH26Unawa
r1Rtf3zLsUtwdJ5VI6au1VjFxeN6+vqwvwkf2N2MsPeQbyKI7/EJjODB3ZjGxSa7FGHUbjblt6j7
S2T7SDpyPEP14QqPx+StNcDkNdRRf/ZIPHmFqKRpXghqwZ8LXb6gggLY/GkG6jI6k3Vu6sU5YTIX
kYNFU8YKr2LunlhtuUfRlpzx2RiJRhPA8Jz9h1bLuhKAl9IUTgVC8joL8euklI1MrOvXQg7rVLrr
v7Rakee9yhkWzI/ACX8gwrZp/gIrSb1xHJByszV4mfwruQL2vvCpOnronkXvDapFwbTCrgoVrm6M
UL826cP9nr3JDqPRhLmu0iMRPwJ6lTHe94vG7IxFLNcf8k1FeqNusBntDZSLxV3gbGj2fCEHA99/
AJ4DdubatHFdlku+hulAsOEwwkvE7qgGnn4pXaMQbWCMSfTzD4UNfdapAlAwbj75tNhbdOgZHTXo
q3JwbGIX/of5XyGJ5fuliA5PDjjlrteFQy1ulRE8NQoWY+clgxQa6v/4gIIqXFpn9codQIZoLg+n
RntB87R92vgW1rRg4EXh7pZzqmLQJOmmPEwt3ZDdkWBbOjyH49YVaZNqpd46kLrSr3X3yvt3YQnO
xqwY9UAWzIRrVLJRLExGcjdfXcHIB/VZZBxI0d24fCw+i7aJg/Z/s0nx5HmIUQ7dctjazjwUOVFU
fJK7jIfPiGRhzgnctyUNtbeoxHGv4Gujk75sa0QSMHPwz8gpQ4XW4k6DxqqWiCGhCElvVSRjpHqX
iOX+i6qCY8/tFStXqlr2twd930+0vlRDdT8KU53645K4is+n0/7smKYWvslGn0Mc+hEvXf45soQp
i66zrIrpv0mggqXQMYykGbSomKP4CFo3ZgRU9FgaxW/ZTGko8W9OD9uQZMv4xhnUCE6vvIIuPypt
aXye30jmr5F0zk/wllSdP0KVo24c+GRouAF5iiTGFn7SlL/DDsBeqm0SzTJgZNqEhdL7BmIIE6vX
ppOT6BUzH1rtv/IyhjTH10RyrqMQsMmxkORGDgCso8VnEJMGtEbSnvASYMpFDfBQNoVU7w5Pm6ha
fXY7RZTkkKshANYrqqdEsirB5yt26yOiMYF38qBgD8w3qrMP9Lmh9Yic+91Izsb1jHE2OjiUmXxk
FsRLVm0JHDJg+aikVXMTPRBXhM/cTmZSyK9nAj9muhbIuwQOW1pXYt+IkB98tu20+nEcqxQvlR6i
yO7DURhOVycF9dhgpOc328UQXIMLDKsYp/r4fidWMMk7TqbGWMm95d4EDBTFwH3gclkc1A4xx2iq
/KOStv67AsiXHtQ25zdg+R55j0qBWckww0XSpBryFxRB0+QVgy1dnKmDaRYk6pW1JwsrQX4olqiD
MtxCptliXt2ygMhvDN0fHAPeeFAa6zHacnnnTmUR+cXCqe+P5UsWynWCyh0N414CmY8O0Q39AWGh
b0cRMFQzQ2BgCknySvBXb147VRHC0I4d318hEJToPXe7SbdUwg12AI09QoSp+iUDaft5E94zUghl
iCscLJXW88zB4qd7Uh20+Fw41VO3lShuRc0wiojiCg3S+pv96xskln4CEJp+fN/USc/tgoDVIwza
CLcJKyImgT3y3N48OBEPvt7lJKgs3+DMAtYfe6ocGb/JoKlIQnhHZdKupjuC6iX0fc/XwADGfezu
IUuZqah7CPffPTsMD+0VrTVxsUFZZ/ACbiyEh9y0cBwfgjimArOZ/H2+YKUEkMI+IyhZTnQymWgT
7Rgj2B5uh94g9ZdCJK1slKA79eCOQuU3V6gQJUpTNvNI96nfdjl05WjZloYl4dwpV0OO0viFnVx0
2Q4QXFJHrEBWOVqDUGPn7iXCZW1MjbuZ+Mnf9Y+7ajQjkzFE7aDewfUegRH1PuYiyuPTe7sMCNxj
XrCX1XGyNgtFs3bwQnU6DS13//L6Ux3EKhqwYr5LGz4kjkrHFS39S+BAiypyX3jCR2NDJf/reGrB
8eplPYbvuTn5hfquDCY3iSHt8nzadIO1a/XY5KaUUgPe9SEeXns4Baw6nZifg12p8yG5OqX6adX0
KvsJymy6g+Z8BG/8E4HYFyoh0jbTMPCHM2MIDeGb+B8QxXDRd4hk5St+dCrCjzJfkj95H0qPaDav
rNsTnl6b8cplfnYbAerWUD9FSmrnRJXntDhFscJ8fxznUvRX1p72rzbjSgOfy+3HTzvaS/iB+o+B
NYk4TD1hm2P6r/EeSRhNLvKtTuD0hOrtIyd2F2U5MDWg3+YTRhWFNBLVM+LWzU6XU+eRRXV5LBwq
MJVvCbVPgIjjwz1cg9CTlzuUFcNG/0/KTJJV02XlmECQt9aDa3nqKBVUHCIJtfl87PHom/3voTZL
BP4qboHgvCrNAJ4RjI2dZkOVEwoDE3UnYQQxMctAlThMYah/u+sTXokinK1Q6OZabS5Wr9W9+DjQ
tOKTXubR7B9KoWI4o1LtUVhKbkIrKUyDj3TRJN5l04KM+pcSuNAW7wSfCHiPYJbTLL78giA9RsCj
SMcRt4hlX2AkTN+F3keWjJY+p5qynXlsQ9oogjgK1mTykOqlNNV9CHeFJmDkAfyppDVgEu1BQ2Yo
gBHuXZRm8L90Oa2VwXYv5ZGrwTO+pf/GhJHSHhMEry/OvVz+3kL+dLkDFil7h4OiENT8D9TQDTen
KMo9ziDqQUYwNDdV1OanxiyIZbwK/3ttfaRS8i0MjGORZrYOo558yL13XjPR2BILspQg699GBxu1
39aSQB2Y0XGu4CW5bTqE/XzLBqKTfnmJK0jiNHyelTHguTsftMGYW7nMTheIPkwUEVIrCjpIgWRp
D7K4i87G/mmcvqtxtoX6mpOxKpWF0kzECYhiUE92OiuD0V4DR7/nAcs5pOOp/OaaOykliuRXkY9J
4xPOkfGRoRUa9sNnRyU7jKxO95prWrlR0tUZ5L9SUwNbknySr4tomlJGznJqDtKnu5nxugb//0Zh
5oPMzAz9vDk2/n6mhK1r0YYiFZXsRImmAavRDfDhlZfhda6+h7CvbYNu8hFlBwN46/eczcSAb3kz
y14L4b+9uJHnkdSsUNhwuZNQLCOgJ4vSqbJ7dNJilWtLzSo4JpCKq27aimF1KINowWwU7T7aaqfz
g1EyYDoR0JhTb5Vwh8/lqUX3y4vImMQF3dXVXppplc8rTDM8VJYcSGfg6YZL0/jneNj2snNZ3VAR
urTqezpNoco+PowKpeyW4mycAlwkg1kMACW1VlLk0eSLhYirZ9zEV7/LsqVm8JJkpk/dklbhfakm
lI/D1B7W3FoKnTDv7FmzQJJZunnD4J/Z2e6KmSGk4TuTVnwgTXNkZGimGjg/0KWeLuHJCZwzPNQE
fR5CbI3hTavtjrkAlWOxK+xp+cF5wThKYLBiST40N0sy3X5T9M6kOffL1/LH3lVFPnQynhGQ/6ip
mL5mFFZPK947TNeJGZr7Mhzb3pVq7PAc7eSM7VABYQZ/GovI8Zd1rEEg5rSn2q3uRcs2teUBYlGh
DhrDPKSRI6aPiX2Xf+6fPDWpVhroXjlpUWWq1yEuDahU/TSD7XqXxMxWigDabtfvGTzkD/ol2yRI
6HaH4dYCo//+wcazA6uIZM0Vnz/rhaExkhG27P9nkabYgmzrHmxCVEHrmQbY8GcMJxkOQXo0Ys7X
Qr6nwC59zUpX8OGZrhMbJ2XD0i3x2ZRXDhO6UD+8BLiX+12Tqt3GIfruwJTMEJP0XhiNFBw8aygY
Ok3cVBuOlQuZhjRLCpE2kIKPEllsYa4G0786uBS0Tv2xGIX3sPZHRq7cE9YL4o0xZUjCDr01UFar
OfKxPTH3mttxAf7wav9ZCVdMRE1gj64xoetR3UlvG8RWeaFQ+nr0S7sGAIU7jG4jn90FTxF5Apbv
5++PH5aA+yXqum/v2fEnFNI3nTXbftwIDfZTH3gnkCS4e93mWLM5apXEs/gaJVVfBH8RMz+PN+y4
zqAja3/K8gLIid+pHxi8ZAt504C2WOXG2FcJxESUd3Ijcxr2e93GywremCGCIHflx9oQuO15IvKf
KJpgGv076mL4WLd0oHB8ZreDdQH1l7q0hc7g5JjdEUGH0u7gsg/2lke8fol2SLasl150napJQy+J
HPP0c0o02Y7BWWoXSx8t8ZBN91CQo/lqU43fXXJhYIFza6kTzksH1vrmv2JFZnnxE3x0asuXEXq2
TA9Wv+ytMWe8c4cmyglGQ+y57cMz9C9FR4kluc8v9wj25e4BpU2k30MqPm7cN8WvvLazE/NYuJnj
mF6UfWgmqkRWx2RfY1rTp+8bB9GihaNVaR9TZAQJoJqrzrHcgvX8k/w8nky/fsDOmwI8OvoJLTWb
nIlWj7JwWA1Lv+KV0Bkg2ARf+zJLxy1Qne8CIySZJBDsZ1rV1rp5QnB4f0HBvsImQL47YC+xhh62
cA2TO2Cfo4vutby52fkyC0h8X0OGlhPdcV10oquATY1B6LEVTqA2F0g5PYaCZkmzTwVb0Caiy4Km
TLCujpNuDK+KhL9ky1vTnstVqlwrNlGpUHofOFbZd8DvaZxUQhxMpaj0AkF6756jIeZ4leUh+d1X
E4oObfpXyK4gQTEsGk2wk9WrHXMcl8NsERApjyXnY6NeJ7oI5+G+oVV3qso9aUk+i4pUHxSQEJif
PRE5/w4U/pZqyWNuB8ZvhYn+PNf2Qhbl76cuU7QQi/HG76fXd5wMVxDNn5vAjIUdIhbIUXRVJLTu
hVDr+8YUFdRWOUxLdl3zmPgEWFkynJM84Utrqv4yo5sg/NKBDdq980UgBv411lL9Y5QpgOi1g6E+
LXMy0bw6VvmihhF1jaPzbLkl+CgB2SXY63I/D5/K2yJvQ/egzH891R5+NcVXkiq37/fKaCrKhHjW
j1vDBSAuOg7XfH+ZTuD7P7iw3Gr+Nl7PYfiqWOmUcC8D5G3hKXSb9Xb5EH8bq8C8Z/+3NOT5a9l0
S/jrvz0I49zVW5iu+WOID4LycTKXFElAhohNbTluqmbjb2p6ks+8hhDIRhM+HJNoCB8TqfKQZqtP
ZMgR/O1urQvoWslA4M9H6XiabeH+TJqmeLW6JQOah3OerkbTwBquy78Axsb9zKdlAL7xqdn+BiUv
l3ZjmHmY2fSH1TWdGJdvMryBIa5/CFwllqIuFgYVEoY/3M/LqacbN8VxVBuos7PmH+htfvDotGjR
Y4Xgp6J4OucSeVc2Y1dMFYLaabJP6KeylBI/bJALVdgt+PbkfjnCV6ZTqLwDVQviKydPuBZVErXT
WGmMpGQrFn/4UXYdT3WPpTHBp8XK/z5kGylm32xIWVpfQp9DBQ3/nl3FLamG00iyR9UOOIgdiUVb
+ObX/O28tGCUW/il7+uDb71lY3gRYWWHwwafCO0v+8a1QNi5tB/F8HrdPhiHzQb2KFFLDVmwFt1r
PXRvDMVrRSMlXgYr5LwVkNc5X2D+W7mFrOKujsuF0puLtZHuMS5vMfh0rPSOrdk2GWmdyskztJ3O
zm45rGv13NKVAaeKvlOytO4Ss4vDNPhTpTF5F+Ssv0RdfmxddQhC6Cks4a0m8D4X8RXY9Cw43GiT
RQgM+GMfYgmolhuEucSqHHSOPb4DcqOkCSpys5K7NEdkgNZh4Xn9QxX7441Pe9AyIO3pes419o6q
olu37ItDCeyslA+ZCDT4dsovo3EHBHlbFSl/je79+21yq6gIG5HFcxj8jWt0Hf5k3HcWMhrnJI+0
ThIxbby0IRJ9Tk+4LcGnM/ZctCWSW0I1HzmVpNKCF38OCXF20Fpmnzs4uVK5PQYjzoxieecX+0e4
u4n8uR8rx3BXuB69gQQb/wLc10kCFjT8pedRdSd87gAsCIUB+cQFrgm8rRY37A6G9VnxEP5Y5lO1
wHrc5vihtrZsTDCsMLRbWQLE+j+5b+U6IuTTryckuLzC/W/9lYFMcpx1Rme2O1KkBIbv0PEYrEgs
LZVUaRhKsa1vlyvQzXNubrEhcJSKcG7U3T6hxRjwsBgnVAeLzdmKPbk32WyZWqkvF45PNoLEfvxX
1+GaIUKOu56MsA/tZ39ddFiuKi6EHhuEdNCUSabcZWi4o9lZJnM6gnuJhC2VvgZC+PFjU83hdj1D
gOYWXPNp5J4aDGGXSYbOBBYapuhSIVK/e54GjJg1MrXbPCCuBDi0PuhECTBXmplMJF1ucciT0cZ8
n54ESGjTif0cTOie6Hbh/CmNQugij+3/3cvspxYgqc3JHanvjfYrQz3nQwZPtC2AKwv0NGyDUzRP
X9YildQ3LiQ97jw3zPEaDWmgxCELV1nKGizAisOxSLKolu3Y8vbxQNacdWDCzPXkxbLMdouhpHnh
lj9FTfLwwDIsLfpg3Jazc56unJarNOtq1eQ6PppOdU3l59Hna9hzFaY+zeJ7g2z7QAsCx9GOEHGv
hxIG83JB5kxA+oMTvo0XYZi9rxSDGyx9Q7w1Jr+3rXae17pckQCZP4/OymPa1wQifA5r/Zq4CPIh
UYrzSZjZa5aGbrlZa47U+/SYWUuNsIiG90OEVABYMdEOwcU7nVaf8qGAexmf54K24NBO8+XCbJ2T
FN90EfbMF/xLrKVfmARK3XivBkBvvW1YecweghdmUpytSjQe7SYdcaQd6Emhi2jOIaUyeha4sW3f
WMReBqboDdMAbeAQsjSY9ksKQRnRPlT8Eo7Wm3OWyEv1u1/LcBLZ7YYSan9gyCmzZsf1cZLARe4s
6hf5fAjhDbOCGa8sMnPXkGJlDw/yDaf+6od5iSRdAq8kW4HrOn2plwTS3tf1Xtk2Mxsy9aSV9P3Q
6yIbrXcYniedV0bzzKO2tTs3bqnOy3dYySa5s1De+NpRRzbt0QDcn7GfP7iP7NA96WpS3jKE9E+g
E0AwOWBJ8FJ9oR1rGejFIPbPziOioK7pw04fIsNgAUiIUwzdzPR7V80pEOr4uwvctE8i+7g/00f8
QmJMK1zIdgOM8s35Bb3uPchODMlsBFTqOKt0jTjXijPNsHhHdTMetyvSztio87WwpJKuhFc873yo
be/acSDKbG9WUd9zRNG6R+tJS2+r7T7i1wCMC5UlLujGvjKWiqTztdxs7363Sn3KSbOjZptAbc8s
3lzBsOzf8oiqeL9YI/dR/zRf4vO1h+EYjHz4HsClR7VAER7NNAurM4QnVZDnOzKFCiSPkrM1zXzc
99LEFjVA55bmXFjAPcSOfH7a4OgDiWhgNd8vWDrMIKAe1Fo/HMXv2xi72V3VGunEkGhPlIvIoJ9U
JZRsFx6EaOY6ooX/fnjLfmkZSv5pdiZjNegrgyM5xkRaDnRkyU0+2rTQtNjkFamBdGEGb3c1OVYA
sO5cieyco+j1QDaw01hVebxYjYnCczf4c4rojlFlfhqdE75pI9N/Czt0RsQfbKY/rwZBFYHKjSSX
ULREYCFHI09/mZBKi0sWcdeONYVm5kL8MvjASuxsHIZRnTKBQpfeTbibTgr4fwhdAHox73jVZqTT
HaZ5Am3lEesfGhz1Dl0c8rG46c2cLwQeIr7+YBsEdJNDkq82pjkE0K6TE7ajFgYIfb5zDvTrbJSl
zmP/EnpNOE9oRnBJrbK1+N+lzcjPH9/6akfQJWnmSCLBo4nVZmK/WBfFIvG5634IV+1HhB5OCt4/
hNG9v2cf9vZNiDTA47xKb/Y18PKJZI9hP7yNmR264+HHIcIUBCtZfge+wtmhyX4RJ1XpyxW4mBeG
IH5MIAzwpVSZDAF/Aiac7s/H6/cIDdc+AZTJ2zwOIR2oCJqTaRFvhoTo8U+EMATrL+a3esE8kvEh
39MQryBhLiz886ZPzeZWmyHseDRWEi+NPvaAoY19BOohW1+cylUQghEbkcFG9ZgHQT2xDvUOLT4S
PwPGh6DDMIZxdsKRxuu8yZvfV7ixQKkw0aQxIvAUHggNPYgtez969uQIzs8qjBGU5l3kgThrQGj8
k+I3IlivRs7rMtDAaOURb2wjUN5BEHE5whjbV7mV8HBGnb5i6JnGGw5G698DeVYPRZkMoePkxtxV
A6tgQ851RgeSn64evqxbkve+GMsRHZUJ8NxL/VbO5xDERM7F0hIKfntlMw0oyZ1lCjAWoIKvt5m7
QD7AJxKxxYm/cav2u8sn4iDlgwZvFr8XoaZ9qKdksPByy/Vs9xWZlrCGBBHUxSLtzTrjz75B7CRl
4trfLeVb6H0LjREq1E0QkJ+CQNMAXnZEo8WObkSuihPoZnldmgiKmCVI6Kh55PS9AjgFasQIftvC
IjX0ueTbY54kn8PhUuz+mYEVzf/ic7U3TauF28BNUu6rR6/KUU8yljqJ4MsHXjbnC5mE+AYg5wNn
Olx4mjCXkgDW4e6UOg8cMFW64XDMmyW0nvJOYplo37T5iN9dJo8IgYbrZWvM0woUoVJxjZqxXWyp
Te9uEoG8PIBd9MEX9r2VXD1zR7JopP3hdab+rL9s/ALfmTlsSOYabWfVGs6y4+kt7F8JHDiodmi9
p2kDiWs0yQGQnHw5quvKz85OFq/UVf5vNVpFlNVFKZ1zi3i3R5Rp7lynDvpskwPGO5DmX2S3ruUA
m7HjgIaBjIzhKRDqzJ7IJQmbLKrFLdaHNezskww6QoVr/hHEY8Eu7nEtyq9lXfuJr09cxTWJHgx6
W1eWBw9B0XEWOpMKcX5q3ajUUMRHhs/JeEwpX2EbOTqHwafmoN/8+ipqTqPzEMlKc3kxAx5zQQQY
cC+vJ1mgSV3FG4eetBQqmk0Qx9r0trEva7uxIMDBMCC+/5mHPG4ffrqUF1agG+KTyze+agjuaT9g
uf7IsSzOlC96Qj21Gxe7akDjJ3R7f4N9szDDJmNgE2XlAtWsWdKWWx3luuEvX9/nt/sckp/MLeSv
KaOEL+FhKQJaFsl6Tw8Y/XaUb1e1TaaQwU7RljYiGaTMLJwvK46JRtq2zRDB/qLNb7+OAQ7lG1hB
i197bEoGv1bY+14cn62qefbk3vXMHMfw0gffrGfH0ZwoO2FLT0tSs35EfDR0/m1mo09M3CAQyiOY
U3QY7tdtprOBDgx2vQ8fIMy2Ag04VumhlmlCOFkwIVfO1Igr900hZzFUFzFZTJpbiuH7J04fElRC
WLlQ1ou8BgRqC9V57wKS4bp00NObWRtM1YtPE3JPKqTsjbC56VN5Oe9mRs2iW8iHeHcNPEbX5dfi
w+SJHm6HnbcBNsk4+o5pkhp2BziWiGy+ZOXrJgowVhrfYpZFXfzLQMrSa64gFTjw8WE3rscodNMb
IKUFFaKXze60SDwHMfZnllNvyWv9YwXWbUk0hgntfqjZu7ZuFzm1UY3eKqaU3fOzTVSWcWeJsVGz
UCNE22IpIfqTVHwyATnlKSWL7Bod8adxSrw4MaBwHYr7lUezxBzgVGaHIv+zy0a2Sk9uXQnT6S3p
/fCHM0Znzp1VW1mDZGB4mfImKzL7FpJWBQd31Rpj51VZS/4wBlyWO4kUz4id1nP/FWk6ctpwScCK
QMJAjxHNPxymigLUwwXqyU8jt7VuxNMAMimxGvb6EnxQBQGQ2MjXc7mGVgMGJcS/8Sew8EHIBYy+
M9/Y/whucW0c4qL6UKocRPzkYYp9jVBprOSRRwM2uhO11Ce3ayR9CiVJr+i5xeTLj9OQPCfon+AW
2fviRoYkg2z1602WB7oFWcsAHs24IqaWADGmjIZVqbOtYKj/c1CrLGFlIiuVOLySKrd0a4beh9Sm
7y6NmmQuKfsCSs7NzaQbIExIrQmPZk9ZlkoN4UKGJRKa+n1F/jBIkyQ22AZvuw6TStRBq+uDWOS8
yO/7T/rQ6GNKjjEFxlYRpeARIbquFBGEOpJC9iwqu8w/f6OVJfATBaqZsyOmx4gKIy57xEZBbJGQ
o6mWAaxqby8S9BkjpXvJYL8d9xGDhtne26t+FMdMAHYfVmDiHk0Qgy7W06oN835ovYUgDQ98IoRl
y4RjKgyBy3FHuA0zF/wSKvpy4Uxn/THbliRZAuZw0BSltoo7G8TdyEVZnngGVxo6uTBlgMIxrdL1
G8frHZgggDrrcQ3mu0Sj+XsD0Kgtri3UpZ7zQbXlaBI6JzF8KpmU4mFmVxZa2Bo1RxBcyDmXJPQ2
qUIHfpcpTdfOOIztJIc7oBfbGXdlPj8OghehnBfnYB7eTJ0hrHoiVZC2ZjsRuAdQNXkY5lDCesmc
pGqMtxDPgCWIdw4WPioJXZ2Yw7cHy/8oQVJQoDGvUcWlZjKRoPfTK/F12UUmt5ePB8zJppKvCZsh
CqWXX4qAXYv+QY38fS9RdbKuiwxxgjA+p8rOa4mhWIlc2sF0nP6l7lBfUvYpO1sia1xPhpWGdKAQ
aaX+vHHrA3/97eDgA6Q1gYvnROE4ER10TYtgU4SUHQS1GIVFMP87vbRT6V59QAXMEh/fTD6Rrf0r
9CIn1xqHJ373YuR5OuND4oebzenLUIlXxxms0s3yUZg1HaWtnRzxa5rkOn7lDzO3gw0J1LVJlE1/
CTZ2EffnYluqT2XcqTc7gvfGIRMprP2jHOgbTZC7b2fAQ4Hzys0p54NKUefPTG8IzlLlq2VJ2+kb
CODAIJDzO5sZQ/NwzBtuDQuSWoOI5Q9oJ234LFk1xLizBSxxcqzi1up5v37bmT07gHFXlvV+UJXr
ksv+nbjB0E9HO96FH08X1jUI8FEnYRPuIbbyUHuLVHd0tCp0TH+2rzV0gnUssV9PhWm8JLwblf1y
952jvmW+MdRnMHLy+EEeJRVktLsIpJwJa5q2+rYYW8R5EQvsQ8/O07WJ2hCZqV4eWHpusU5mCAJw
v+tiiMWNwJNZzmrs7edefVh88P9fm3gWrWaE/KcdDJDF73iExnFEeErV7/Q589Kfdg7WYPl0M3Zx
sCCRmnG36+3/831yxO4ZBfajpZWZImrdA4mNjzQdD/Vky2eqOysHa9X05PUBN9nkhhptPOfo6lqu
6DNRPQla6RzLp8rjLAFKOXMnVGfiCWGm2LHrvAocO9xMWCDa4sGSN1cOkiT/e0lfzJJ0VJh8VGjc
mR2fH5EfrMV2F83gdqLsf6Exs+7leGDnFAodPPJEPpzdnx3eOaHC5V13ScwxIUVQZEtL7VVJ59Qj
ygS5rIiQEDOW3q7k/bxEQuZMOtTyczQgXK/ejCxBoS3kHRp8I7D7YCaSqaYepSLc0mi/SgUYBlA0
25A3W1RsnIEAOA06oq3GI6tRY0r66A7lmvDOainp8uIFGF2v4t3LNL+YBYyVmEc/bFY2Y8mHGNa4
LldL0QzdkpcU3I7oze/+CGCxGz8hPk4Q7YqqRblLMPoUbR4+A/XJ7dOZ00OKa+3WPYdbb1K7aXbM
2HDDWJ8HyL9jtQ36QmOJvaZo/TK8swuEVpsgKbF0hj441XpNcw5f1RsIX00GXqAM7eRglCjpwQgE
hfFVa9No/WhxybmRM9QyeiikNMyBHX3rRvZzw8z0wJsT8atiOeEc3G3GWNkXtI63A2AsA2Zwe10u
lB51TN8rksP0UrzS00vcddQbQWdRrxqk87/oNape8Vwtmzyt2YC6gH8EpO3cqR6RLNtB81EUwzMl
UwUu5FtdIzxjLByRJWvDenSC8rugr6FYo8N4mQqmvAzRFDvfu4BwMqjohd4812536w5ayc0Wj62h
QXV1JWaxwKh/NHG1oH9JL2ctSZQTMxLRld/QFn2JaP7YRuFE91EPES2MFPfngQ2fqBJMoDUb/ZsG
dMW9ccqSJMwlBTee67HJlezVBFAcjjDdhgubD8iw3DpmGHZgegFdMrspSaCjWFSGDpnB9/sYO5VV
DEdvzclk01i+zNH3myZtc4ykiO99kFS+vwKUR6SX4hO/WIK+hJfXj5Tf0bZxecz6xSlmnT5FTQ99
or8U2xLe73lAU48SFs2gkVEVqcnjDPL3AV1ZdP1vrW3TE8T+J9uwtHjmtES2uyy252zLzihE+95y
eF5aXwomCxOE4bqwQjChtCbkudf6cwP8pJ3zuRvxMpG9Jn/hkFIL5FqU0lbEbZY02kE9iaXfQxFZ
5zQgcKMDkbLmMhPLlWmFAopqnVQQRKDjxpQvyVSfU/U+NxazZzCznjfbZp5L/hfCgjeRq7LGnbiA
T5j7Jw7q3Xw81ez76VcZBnGE1CGvz/7qDg7Fl4nUzWBwot+mrPNq+Ky55nxAD0iKkWrCUP2DgyaZ
EGtmghpBo1Fau0g9/rhA2v1hkJtDAnsCaNkN3PZpSYEzto9ok6S3pBc4uCKoEn4Ztj1BPsnQKlqs
HRhBd4zyK1d7XVgVrlG4Vj37DXLUaYAvYvfxk3lMjmioUFjBwK+NtnRjXtyqN7SxdiyOdkMTmrBF
w3VEDJANCuabbJm/uYKFcbm8zA7EXmQ4iMTTgR37bLPZaPFvTGJldFRD/adVi/OYIZ2C8Xm55KpY
kVvgX85qY6jRTsYo8TRUxNr4PLQ7+9wuvCCeynAQWB1uxMlwHLCKKrT9eod4tIyRUMkGQrA0t8qs
Gzo98nnytZx3TnXam/qZ3VWlaz+VWk/zhcTmqezflwW3N3qPsXyr/+L8v3PWb5Se+K9hp/26fw8S
TNPHbp4IsOh1Bls1/wLxi6GYQdvzVaMd56PAaqWHLbvhKbMJLvlQW60M7/K1CHVDC2DQ6nMVoV/p
2N6S219BDsd0jhIlpgngig6qpNeXgIR8wCSq094YjeCmOGMs7m4VaTI96VfVNWR2CZ2p54KR+GUT
YcX1qh6d1muQo0FFDiLhwBg08f47HUpLZihEf6JvGcHIYsXDu+ss2gSZiCz3r7zh3cJcKn8ZMmT9
TUIxi55cp6JBaY1R8HcjNBVgRoGiXuPJxs+9UIPujemtVsH2328ErVYKKhSybsuM3KNNR9G7Rjee
El4F8bZMSxBXHD0i3uhilUpMf0eWIItwOCA4hb3D3qncwtVXvdBe1fMUfbpkP2oZrx4hZ6FF27vu
SZ1UEB8A7hn4fA3modnhbNysuBp7IutFuOqHAxPtyLmiVPrSN01aMSRVkJ1G5OrmpuN3FJJopHHJ
CjOj3cQe1LIpHZiUbxaMp46eAtGIyROukugtfTff8kcgluQ6VUwHkN5RcarG4IP5bqVyA5xtJKcY
5MTSacJiR5CirAs9FEhiDrNkQaqrTQli947vRct4Nm+yaqxSFBEsC3hkuey6J6wt2Xb7hLmRX0Ov
IToZuyrgB3TrAIffinEti2wuER+kk6K2ta+n7S6YRAYguff0TXaLKrqXippdanvr2Tk02sadMAWt
z06K9cra79xk4hko0cl9bVsOjVdf0se+EcqazJ/iVsSZVB/uLARaPTj5+pqAW565t9IBKt1uZQ3Q
AGCIL+v5lJWN1ZuZopvNaei6zT44sS6sDwbrIxqLH455ehhhGsgUeRzIrkPGtmW7qFpy93nxUQwb
UHzU3Is2Di0nPgYjnV9dPbHGm1MNLMl77Zzhpn5wDXpIp4Mzpw/7M96Gedi4EieCAwoID3AE2iHc
liy8RP8ltEi7vRk0ElodFHH9im/LmylLqlcnnZ7sqESljdMYbbfcRsefUZNMZsZ6ZrB+uvj8PjZH
+hegdX45OWxQS3CX0iD4HR66pOrULboG2855w1P43cl+3luqKGEeIJoK0Ytl8dXxc+CX0x+QiSlG
8ZL/b349S5ZJQLz3V6iHMHmb/gNoeypdCJc2h5WJMcgZu+dEd7hfoeqY9vyFCXZYQZJU4MVV2Gg+
A/o/X7EwL+TZTmzSOxVVIC5M3IR63B1yj10ewtJcivVoO2uKvs2FSZCAWQ1Ghb9j4ggPxVqpPZ6k
Fx/9yBNYMiXULy5BO/nBAUs+hayZKx4HSNq170mPffYRxIoxLIrlm8bBYpSraXljFXJ/Ievo4/wZ
AgEopcAnAiPt9yJ9odKap1cFhQIdc1IzXUu73QgTTz0bClt2a8iK+mxNgiR9h3+/RSh8r7ChdC4W
5yoPCUOsPojc+WcwxsIqkhWqK+g7ZzaMDJbVSOo0PzhjMQRNehXExKQzm6YvEccgSSAnUNo1LQjg
d5EG/r6VY0Sk6b6Cvrti7cV0J8BPHCWxJ2rYnu9NYmbtgT4KP+p/PLjECI0weaQaoiv0Hn/ai5hL
ONeqC2b0/8UiGXyd/usvcdwuieEWozfdaBqv3gn9STaBe1g0JiHfJGHJ55VdnyRljYjwfRk/504F
U7nbRZus+KoOGZbAD5C9+F2vFZedop/o7+H7XBjpaTK8ARTzeZPkf/tCkL+FkXzIzVkB7I96UnUC
h9N8SBXfZWYxGHYZKvw1/s7p+PBHLo6vPnDgVynoOkOaoD/Meya1xIFQTe0WSsNO9LCtXJVhaPhd
iXPG5YOc8Le4gH+TzUnKzWtoJbag9crncYrP2MRp+YluCf5DFRZCpx2dfld6sRhdEmrlzbbJYs1U
F/mj1lFG6v+cbvjdxsajL+Dd6/7+FFBuxTVGe585HNRtNML4tBq7jgTpsde71GzjmSSxTb4AVVvM
vLITVbHieGmE1STr3BsekGD7yHe7XTK1/XJOinD8NhusZFPOKTp657rWBnAVjxVcHmEquo4LhBNx
Y+wt55eAeE+0UY2GOCPEZmsb/IyG92LI0szn2m+6ZnsArqddhizGhEFpkaRRXIEWea3Z1y11JMRA
4TeFYMh4jFW4D6DeSGFauywhUHC6WPG0Xnl/Xz9EWMDBQz49Znq0C1CHkTwqk1VWMMri5uXrdLS3
59g7D1pEe7TqVjpVXPw/ejC+JszMP/FtgCla6StCull6lEKU7lRKs8Cmh9TnnwqZGslrVvSLzxkf
8ZQeRfHNZEO/drJGdzeZainWVbbJZHWg4xSq/XxOHjTtPqepJgkCfg56AYHn/NRzQ5gNvmVMo/B3
un96OeGYW3pFRbkpYRw4XNlPnWzfwb/OVIR042uMGzqdufKKUlhk29XOdbegqEcFEZ/iBRUGe1oc
orS57aMQ6wlfZnCP3VoSG7t9U6+hKmW8mrXp2Gh3pSyBQfmXMhp8pSE9qN08TloYHnDalVYOYC2n
J0uka+1U3eB8yhKJ5uMNAh2h7qfbsFVybl21mynDrS/6OK8JWGrOP2al6S7XriyK8cBuEx5WcO+X
Oq7PJJPe/5UHp/LSDl5XosNqr4SNMqKa39vIn3+9DarkFG3f2fy7mi6muQO/C9dq0k1n/baJ+taR
mkMlWR9dtjJP1Fshyhrkj5lLLJN6xHTRAJ88egUQyBIfLnrIf2L7dsLdjIaw/snxq3fqMzwCP3Yx
MclzXWBc4WVbZ8QlmCkScMjh29gwbNvhs46Lza6yuo+XWaU8Z406XCDlQ3IVuXiYbUH07SJZTpO6
G3w2WWPmJT2eKMbZkRiw5qsaVcukPYL/5wkIQgFxSCGQGe3rewiTGmoZQ4PA+XWD7dQExCgIGxG6
pUwYhYCDT47aj0BeEr9xO9bPSF3VHLwdCmsHDVKzexmOHnPaFIVtPYRsSh3pRKNe3MM1grZYj0Xs
EvGDk3fUukI7RglGYYnVe7W04NaY3luM5/MYDXvbiMtfdhcPrwXg7mrgRYHRFSqTupC3gcsZe/Mb
TczWBgnA7GFLBX9jzu/L36IQRw/ZpisdV0ZW8NmkbzeewhF2Mio0J5pWHjndhuYJFqSN4HwPMH+B
FpLMXueBcn4AGBNXq/1wrmq6/9sPGeFPBE4KzxZ+HgON4sllOvzMZXb5Hhs0Ff336J9RI8OXuOsj
CP66lGkc+atOF0QrddOxdTLCaQkw/Ii/YHJdRkfYG2FrwJjK8cYbDJrGm1Iya2t5ajCNBpEC7L99
cA3VMxWNh8KyEPXx8qIsKPFYeOiZaJEmXgWAcq/jnx3PVOMqBhvtd2/asfYfhfFO7nTqavqqsAEL
BlBG5l/Olo9mcR0H5aEMmkDemh21Vp1DCMQJXiPeJC0YBgQ9B22r3sbe8t1WLcfperjHt4lSuuyN
DSMla6XiIIsjfYKkGzuc27qEgQMEDtERR9a4H+zHi6CrhJZzuLPsEUvUZ0vvV+7y5z3ewak9zmgX
e2qflZdu6G1VJg0jBoF8YO762iCZSX1SSYY5bq/JlSHo09WhOFoM6A3zvhlru2gfGi0w7RoRCma/
jNuWTrqMtIxKDf2czWCasTpi7WLDBeB5bQIw/1fVofLBO0hbiqr4Suj2WB6MvikceDhu97NI+feb
Ra9UZQ/+QRgsS9sni2z9xMqNf+DkX1XSD1jgd+JbXMCnlcR2D2VbMry5BThMDrnU12/HFin3HxPw
IXorIEiwk23mBEE8hU81nE/t7nBGTf3VwehKFttLKfLoxuHxkNsqwCz1wRtKqld2ao3/qfHv7PRr
IVySnUYMsGih1XPNtpsITcQ3QVeLboSGxcaat56Ui8AUvxI+vRB5SLI5JBZwJ3SiSPN60RZap5Lu
vuMgia5LgvQhXIGdcFIf3FLOjsHcfOxCe33HRv5gZAL3atbq318/a97rc3iUi6aK8F6Msdbh1uXQ
IKbhZB8rlClut6EzHfJKBfy+98FojaZhxJaRWmKdi1lIN3wzZkW7zKa41JEi9HPRQtUNHl5H8V4x
ZTTMO6t/c+YBDO9/eyETg76wpQVwxms1hLu/buY58x9HmWRsA1kY1GzaJ8ubiifZU3VjOZpGaXQH
kEA1gN4WqTBFUxk/6P5PgpaofHi/6FoPUFHzVYfVAIEeocHlrvxxn+IJ6HOozzAnXxkv/SHDPSqm
IdXZ6iepo2eg7klNsQ==
`protect end_protected

